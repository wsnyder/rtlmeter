// Modified by Princeton University on June 9th, 2015
// ========== Copyright Header Begin ==========================================
//
// OpenSPARC T1 Processor File: ciop_iob.v
// Copyright (c) 2006 Sun Microsystems, Inc.  All Rights Reserved.
// DO NOT ALTER OR REMOVE COPYRIGHT NOTICES.
//
// The above named program is free software; you can redistribute it and/or
// modify it under the terms of the GNU General Public
// License version 2 as published by the Free Software Foundation.
//
// The above named program is distributed in the hope that it will be
// useful, but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
// General Public License for more details.
//
// You should have received a copy of the GNU General Public
// License along with this work; if not, write to the Free Software
// Foundation, Inc., 51 Franklin St, Fifth Floor, Boston, MA 02110-1301, USA.
//
// ========== Copyright Header End ============================================
`timescale 1ps/1ps
`include "define.tmp.h"
`include "cross_module.tmp.h"

// /home/gl/work/openpiton/piton/verif/env/manycore/devices_ariane.xml


module ciop_fake_iob(
    input clk,
    input rst_n,

    output reg noc_out_val,
    input noc_out_rdy,
    output reg [`NOC_DATA_WIDTH-1:0] noc_out_data
,
   input                spc0_inst_done,
   input [63:0]         pc_w0

,
   input                spc1_inst_done,
   input [63:0]         pc_w1

,
   input                spc2_inst_done,
   input [63:0]         pc_w2

,
   input                spc3_inst_done,
   input [63:0]         pc_w3

,
   input                spc4_inst_done,
   input [63:0]         pc_w4

,
   input                spc5_inst_done,
   input [63:0]         pc_w5

,
   input                spc6_inst_done,
   input [63:0]         pc_w6

,
   input                spc7_inst_done,
   input [63:0]         pc_w7

,
   input                spc8_inst_done,
   input [63:0]         pc_w8

,
   input                spc9_inst_done,
   input [63:0]         pc_w9

,
   input                spc10_inst_done,
   input [63:0]         pc_w10

,
   input                spc11_inst_done,
   input [63:0]         pc_w11

,
   input                spc12_inst_done,
   input [63:0]         pc_w12

,
   input                spc13_inst_done,
   input [63:0]         pc_w13

,
   input                spc14_inst_done,
   input [63:0]         pc_w14

,
   input                spc15_inst_done,
   input [63:0]         pc_w15

,
   input                spc16_inst_done,
   input [63:0]         pc_w16

,
   input                spc17_inst_done,
   input [63:0]         pc_w17

,
   input                spc18_inst_done,
   input [63:0]         pc_w18

,
   input                spc19_inst_done,
   input [63:0]         pc_w19

,
   input                spc20_inst_done,
   input [63:0]         pc_w20

,
   input                spc21_inst_done,
   input [63:0]         pc_w21

,
   input                spc22_inst_done,
   input [63:0]         pc_w22

,
   input                spc23_inst_done,
   input [63:0]         pc_w23

,
   input                spc24_inst_done,
   input [63:0]         pc_w24

,
   input                spc25_inst_done,
   input [63:0]         pc_w25

,
   input                spc26_inst_done,
   input [63:0]         pc_w26

,
   input                spc27_inst_done,
   input [63:0]         pc_w27

,
   input                spc28_inst_done,
   input [63:0]         pc_w28

,
   input                spc29_inst_done,
   input [63:0]         pc_w29

,
   input                spc30_inst_done,
   input [63:0]         pc_w30

,
   input                spc31_inst_done,
   input [63:0]         pc_w31

,
   input                spc32_inst_done,
   input [63:0]         pc_w32

,
   input                spc33_inst_done,
   input [63:0]         pc_w33

,
   input                spc34_inst_done,
   input [63:0]         pc_w34

,
   input                spc35_inst_done,
   input [63:0]         pc_w35

,
   input                spc36_inst_done,
   input [63:0]         pc_w36

,
   input                spc37_inst_done,
   input [63:0]         pc_w37

,
   input                spc38_inst_done,
   input [63:0]         pc_w38

,
   input                spc39_inst_done,
   input [63:0]         pc_w39

,
   input                spc40_inst_done,
   input [63:0]         pc_w40

,
   input                spc41_inst_done,
   input [63:0]         pc_w41

,
   input                spc42_inst_done,
   input [63:0]         pc_w42

,
   input                spc43_inst_done,
   input [63:0]         pc_w43

,
   input                spc44_inst_done,
   input [63:0]         pc_w44

,
   input                spc45_inst_done,
   input [63:0]         pc_w45

,
   input                spc46_inst_done,
   input [63:0]         pc_w46

,
   input                spc47_inst_done,
   input [63:0]         pc_w47

,
   input                spc48_inst_done,
   input [63:0]         pc_w48

,
   input                spc49_inst_done,
   input [63:0]         pc_w49

,
   input                spc50_inst_done,
   input [63:0]         pc_w50

,
   input                spc51_inst_done,
   input [63:0]         pc_w51

,
   input                spc52_inst_done,
   input [63:0]         pc_w52

,
   input                spc53_inst_done,
   input [63:0]         pc_w53

,
   input                spc54_inst_done,
   input [63:0]         pc_w54

,
   input                spc55_inst_done,
   input [63:0]         pc_w55

,
   input                spc56_inst_done,
   input [63:0]         pc_w56

,
   input                spc57_inst_done,
   input [63:0]         pc_w57

,
   input                spc58_inst_done,
   input [63:0]         pc_w58

,
   input                spc59_inst_done,
   input [63:0]         pc_w59

,
   input                spc60_inst_done,
   input [63:0]         pc_w60

,
   input                spc61_inst_done,
   input [63:0]         pc_w61

,
   input                spc62_inst_done,
   input [63:0]         pc_w62

,
   input                spc63_inst_done,
   input [63:0]         pc_w63

,
   input                spc64_inst_done,
   input [63:0]         pc_w64

,
   input                spc65_inst_done,
   input [63:0]         pc_w65

,
   input                spc66_inst_done,
   input [63:0]         pc_w66

,
   input                spc67_inst_done,
   input [63:0]         pc_w67

,
   input                spc68_inst_done,
   input [63:0]         pc_w68

,
   input                spc69_inst_done,
   input [63:0]         pc_w69

,
   input                spc70_inst_done,
   input [63:0]         pc_w70

,
   input                spc71_inst_done,
   input [63:0]         pc_w71

,
   input                spc72_inst_done,
   input [63:0]         pc_w72

,
   input                spc73_inst_done,
   input [63:0]         pc_w73

,
   input                spc74_inst_done,
   input [63:0]         pc_w74

,
   input                spc75_inst_done,
   input [63:0]         pc_w75

,
   input                spc76_inst_done,
   input [63:0]         pc_w76

,
   input                spc77_inst_done,
   input [63:0]         pc_w77

,
   input                spc78_inst_done,
   input [63:0]         pc_w78

,
   input                spc79_inst_done,
   input [63:0]         pc_w79

,
   input                spc80_inst_done,
   input [63:0]         pc_w80

,
   input                spc81_inst_done,
   input [63:0]         pc_w81

,
   input                spc82_inst_done,
   input [63:0]         pc_w82

,
   input                spc83_inst_done,
   input [63:0]         pc_w83

,
   input                spc84_inst_done,
   input [63:0]         pc_w84

,
   input                spc85_inst_done,
   input [63:0]         pc_w85

,
   input                spc86_inst_done,
   input [63:0]         pc_w86

,
   input                spc87_inst_done,
   input [63:0]         pc_w87

,
   input                spc88_inst_done,
   input [63:0]         pc_w88

,
   input                spc89_inst_done,
   input [63:0]         pc_w89

,
   input                spc90_inst_done,
   input [63:0]         pc_w90

,
   input                spc91_inst_done,
   input [63:0]         pc_w91

,
   input                spc92_inst_done,
   input [63:0]         pc_w92

,
   input                spc93_inst_done,
   input [63:0]         pc_w93

,
   input                spc94_inst_done,
   input [63:0]         pc_w94

,
   input                spc95_inst_done,
   input [63:0]         pc_w95

,
   input                spc96_inst_done,
   input [63:0]         pc_w96

,
   input                spc97_inst_done,
   input [63:0]         pc_w97

,
   input                spc98_inst_done,
   input [63:0]         pc_w98

,
   input                spc99_inst_done,
   input [63:0]         pc_w99

,
   input                spc100_inst_done,
   input [63:0]         pc_w100

,
   input                spc101_inst_done,
   input [63:0]         pc_w101

,
   input                spc102_inst_done,
   input [63:0]         pc_w102

,
   input                spc103_inst_done,
   input [63:0]         pc_w103

,
   input                spc104_inst_done,
   input [63:0]         pc_w104

,
   input                spc105_inst_done,
   input [63:0]         pc_w105

,
   input                spc106_inst_done,
   input [63:0]         pc_w106

,
   input                spc107_inst_done,
   input [63:0]         pc_w107

,
   input                spc108_inst_done,
   input [63:0]         pc_w108

,
   input                spc109_inst_done,
   input [63:0]         pc_w109

,
   input                spc110_inst_done,
   input [63:0]         pc_w110

,
   input                spc111_inst_done,
   input [63:0]         pc_w111

,
   input                spc112_inst_done,
   input [63:0]         pc_w112

,
   input                spc113_inst_done,
   input [63:0]         pc_w113

,
   input                spc114_inst_done,
   input [63:0]         pc_w114

,
   input                spc115_inst_done,
   input [63:0]         pc_w115

,
   input                spc116_inst_done,
   input [63:0]         pc_w116

,
   input                spc117_inst_done,
   input [63:0]         pc_w117

,
   input                spc118_inst_done,
   input [63:0]         pc_w118

,
   input                spc119_inst_done,
   input [63:0]         pc_w119

,
   input                spc120_inst_done,
   input [63:0]         pc_w120

,
   input                spc121_inst_done,
   input [63:0]         pc_w121

,
   input                spc122_inst_done,
   input [63:0]         pc_w122

,
   input                spc123_inst_done,
   input [63:0]         pc_w123

,
   input                spc124_inst_done,
   input [63:0]         pc_w124

,
   input                spc125_inst_done,
   input [63:0]         pc_w125

,
   input                spc126_inst_done,
   input [63:0]         pc_w126

,
   input                spc127_inst_done,
   input [63:0]         pc_w127

,
   input                spc128_inst_done,
   input [63:0]         pc_w128

,
   input                spc129_inst_done,
   input [63:0]         pc_w129

,
   input                spc130_inst_done,
   input [63:0]         pc_w130

,
   input                spc131_inst_done,
   input [63:0]         pc_w131

,
   input                spc132_inst_done,
   input [63:0]         pc_w132

,
   input                spc133_inst_done,
   input [63:0]         pc_w133

,
   input                spc134_inst_done,
   input [63:0]         pc_w134

,
   input                spc135_inst_done,
   input [63:0]         pc_w135

,
   input                spc136_inst_done,
   input [63:0]         pc_w136

,
   input                spc137_inst_done,
   input [63:0]         pc_w137

,
   input                spc138_inst_done,
   input [63:0]         pc_w138

,
   input                spc139_inst_done,
   input [63:0]         pc_w139

,
   input                spc140_inst_done,
   input [63:0]         pc_w140

,
   input                spc141_inst_done,
   input [63:0]         pc_w141

,
   input                spc142_inst_done,
   input [63:0]         pc_w142

,
   input                spc143_inst_done,
   input [63:0]         pc_w143

,
   input                spc144_inst_done,
   input [63:0]         pc_w144

,
   input                spc145_inst_done,
   input [63:0]         pc_w145

,
   input                spc146_inst_done,
   input [63:0]         pc_w146

,
   input                spc147_inst_done,
   input [63:0]         pc_w147

,
   input                spc148_inst_done,
   input [63:0]         pc_w148

,
   input                spc149_inst_done,
   input [63:0]         pc_w149

,
   input                spc150_inst_done,
   input [63:0]         pc_w150

,
   input                spc151_inst_done,
   input [63:0]         pc_w151

,
   input                spc152_inst_done,
   input [63:0]         pc_w152

,
   input                spc153_inst_done,
   input [63:0]         pc_w153

,
   input                spc154_inst_done,
   input [63:0]         pc_w154

,
   input                spc155_inst_done,
   input [63:0]         pc_w155

,
   input                spc156_inst_done,
   input [63:0]         pc_w156

,
   input                spc157_inst_done,
   input [63:0]         pc_w157

,
   input                spc158_inst_done,
   input [63:0]         pc_w158

,
   input                spc159_inst_done,
   input [63:0]         pc_w159

,
   input                spc160_inst_done,
   input [63:0]         pc_w160

,
   input                spc161_inst_done,
   input [63:0]         pc_w161

,
   input                spc162_inst_done,
   input [63:0]         pc_w162

,
   input                spc163_inst_done,
   input [63:0]         pc_w163

,
   input                spc164_inst_done,
   input [63:0]         pc_w164

,
   input                spc165_inst_done,
   input [63:0]         pc_w165

,
   input                spc166_inst_done,
   input [63:0]         pc_w166

,
   input                spc167_inst_done,
   input [63:0]         pc_w167

,
   input                spc168_inst_done,
   input [63:0]         pc_w168

,
   input                spc169_inst_done,
   input [63:0]         pc_w169

,
   input                spc170_inst_done,
   input [63:0]         pc_w170

,
   input                spc171_inst_done,
   input [63:0]         pc_w171

,
   input                spc172_inst_done,
   input [63:0]         pc_w172

,
   input                spc173_inst_done,
   input [63:0]         pc_w173

,
   input                spc174_inst_done,
   input [63:0]         pc_w174

,
   input                spc175_inst_done,
   input [63:0]         pc_w175

,
   input                spc176_inst_done,
   input [63:0]         pc_w176

,
   input                spc177_inst_done,
   input [63:0]         pc_w177

,
   input                spc178_inst_done,
   input [63:0]         pc_w178

,
   input                spc179_inst_done,
   input [63:0]         pc_w179

,
   input                spc180_inst_done,
   input [63:0]         pc_w180

,
   input                spc181_inst_done,
   input [63:0]         pc_w181

,
   input                spc182_inst_done,
   input [63:0]         pc_w182

,
   input                spc183_inst_done,
   input [63:0]         pc_w183

,
   input                spc184_inst_done,
   input [63:0]         pc_w184

,
   input                spc185_inst_done,
   input [63:0]         pc_w185

,
   input                spc186_inst_done,
   input [63:0]         pc_w186

,
   input                spc187_inst_done,
   input [63:0]         pc_w187

,
   input                spc188_inst_done,
   input [63:0]         pc_w188

,
   input                spc189_inst_done,
   input [63:0]         pc_w189

,
   input                spc190_inst_done,
   input [63:0]         pc_w190

,
   input                spc191_inst_done,
   input [63:0]         pc_w191

,
   input                spc192_inst_done,
   input [63:0]         pc_w192

,
   input                spc193_inst_done,
   input [63:0]         pc_w193

,
   input                spc194_inst_done,
   input [63:0]         pc_w194

,
   input                spc195_inst_done,
   input [63:0]         pc_w195

,
   input                spc196_inst_done,
   input [63:0]         pc_w196

,
   input                spc197_inst_done,
   input [63:0]         pc_w197

,
   input                spc198_inst_done,
   input [63:0]         pc_w198

,
   input                spc199_inst_done,
   input [63:0]         pc_w199

,
   input                spc200_inst_done,
   input [63:0]         pc_w200

,
   input                spc201_inst_done,
   input [63:0]         pc_w201

,
   input                spc202_inst_done,
   input [63:0]         pc_w202

,
   input                spc203_inst_done,
   input [63:0]         pc_w203

,
   input                spc204_inst_done,
   input [63:0]         pc_w204

,
   input                spc205_inst_done,
   input [63:0]         pc_w205

,
   input                spc206_inst_done,
   input [63:0]         pc_w206

,
   input                spc207_inst_done,
   input [63:0]         pc_w207

,
   input                spc208_inst_done,
   input [63:0]         pc_w208

,
   input                spc209_inst_done,
   input [63:0]         pc_w209

,
   input                spc210_inst_done,
   input [63:0]         pc_w210

,
   input                spc211_inst_done,
   input [63:0]         pc_w211

,
   input                spc212_inst_done,
   input [63:0]         pc_w212

,
   input                spc213_inst_done,
   input [63:0]         pc_w213

,
   input                spc214_inst_done,
   input [63:0]         pc_w214

,
   input                spc215_inst_done,
   input [63:0]         pc_w215

,
   input                spc216_inst_done,
   input [63:0]         pc_w216

,
   input                spc217_inst_done,
   input [63:0]         pc_w217

,
   input                spc218_inst_done,
   input [63:0]         pc_w218

,
   input                spc219_inst_done,
   input [63:0]         pc_w219

,
   input                spc220_inst_done,
   input [63:0]         pc_w220

,
   input                spc221_inst_done,
   input [63:0]         pc_w221

,
   input                spc222_inst_done,
   input [63:0]         pc_w222

,
   input                spc223_inst_done,
   input [63:0]         pc_w223

,
   input                spc224_inst_done,
   input [63:0]         pc_w224

,
   input                spc225_inst_done,
   input [63:0]         pc_w225

,
   input                spc226_inst_done,
   input [63:0]         pc_w226

,
   input                spc227_inst_done,
   input [63:0]         pc_w227

,
   input                spc228_inst_done,
   input [63:0]         pc_w228

,
   input                spc229_inst_done,
   input [63:0]         pc_w229

,
   input                spc230_inst_done,
   input [63:0]         pc_w230

,
   input                spc231_inst_done,
   input [63:0]         pc_w231

,
   input                spc232_inst_done,
   input [63:0]         pc_w232

,
   input                spc233_inst_done,
   input [63:0]         pc_w233

,
   input                spc234_inst_done,
   input [63:0]         pc_w234

,
   input                spc235_inst_done,
   input [63:0]         pc_w235

,
   input                spc236_inst_done,
   input [63:0]         pc_w236

,
   input                spc237_inst_done,
   input [63:0]         pc_w237

,
   input                spc238_inst_done,
   input [63:0]         pc_w238

,
   input                spc239_inst_done,
   input [63:0]         pc_w239

,
   input                spc240_inst_done,
   input [63:0]         pc_w240

,
   input                spc241_inst_done,
   input [63:0]         pc_w241

,
   input                spc242_inst_done,
   input [63:0]         pc_w242

,
   input                spc243_inst_done,
   input [63:0]         pc_w243

,
   input                spc244_inst_done,
   input [63:0]         pc_w244

,
   input                spc245_inst_done,
   input [63:0]         pc_w245

,
   input                spc246_inst_done,
   input [63:0]         pc_w246

,
   input                spc247_inst_done,
   input [63:0]         pc_w247

,
   input                spc248_inst_done,
   input [63:0]         pc_w248

,
   input                spc249_inst_done,
   input [63:0]         pc_w249

,
   input                spc250_inst_done,
   input [63:0]         pc_w250

,
   input                spc251_inst_done,
   input [63:0]         pc_w251

,
   input                spc252_inst_done,
   input [63:0]         pc_w252

,
   input                spc253_inst_done,
   input [63:0]         pc_w253

,
   input                spc254_inst_done,
   input [63:0]         pc_w254

,
   input                spc255_inst_done,
   input [63:0]         pc_w255

,
   input                spc256_inst_done,
   input [63:0]         pc_w256

,
   input                spc257_inst_done,
   input [63:0]         pc_w257

,
   input                spc258_inst_done,
   input [63:0]         pc_w258

,
   input                spc259_inst_done,
   input [63:0]         pc_w259

,
   input                spc260_inst_done,
   input [63:0]         pc_w260

,
   input                spc261_inst_done,
   input [63:0]         pc_w261

,
   input                spc262_inst_done,
   input [63:0]         pc_w262

,
   input                spc263_inst_done,
   input [63:0]         pc_w263

,
   input                spc264_inst_done,
   input [63:0]         pc_w264

,
   input                spc265_inst_done,
   input [63:0]         pc_w265

,
   input                spc266_inst_done,
   input [63:0]         pc_w266

,
   input                spc267_inst_done,
   input [63:0]         pc_w267

,
   input                spc268_inst_done,
   input [63:0]         pc_w268

,
   input                spc269_inst_done,
   input [63:0]         pc_w269

,
   input                spc270_inst_done,
   input [63:0]         pc_w270

,
   input                spc271_inst_done,
   input [63:0]         pc_w271

,
   input                spc272_inst_done,
   input [63:0]         pc_w272

,
   input                spc273_inst_done,
   input [63:0]         pc_w273

,
   input                spc274_inst_done,
   input [63:0]         pc_w274

,
   input                spc275_inst_done,
   input [63:0]         pc_w275

,
   input                spc276_inst_done,
   input [63:0]         pc_w276

,
   input                spc277_inst_done,
   input [63:0]         pc_w277

,
   input                spc278_inst_done,
   input [63:0]         pc_w278

,
   input                spc279_inst_done,
   input [63:0]         pc_w279

,
   input                spc280_inst_done,
   input [63:0]         pc_w280

,
   input                spc281_inst_done,
   input [63:0]         pc_w281

,
   input                spc282_inst_done,
   input [63:0]         pc_w282

,
   input                spc283_inst_done,
   input [63:0]         pc_w283

,
   input                spc284_inst_done,
   input [63:0]         pc_w284

,
   input                spc285_inst_done,
   input [63:0]         pc_w285

,
   input                spc286_inst_done,
   input [63:0]         pc_w286

,
   input                spc287_inst_done,
   input [63:0]         pc_w287

,
   input                spc288_inst_done,
   input [63:0]         pc_w288

,
   input                spc289_inst_done,
   input [63:0]         pc_w289

,
   input                spc290_inst_done,
   input [63:0]         pc_w290

,
   input                spc291_inst_done,
   input [63:0]         pc_w291

,
   input                spc292_inst_done,
   input [63:0]         pc_w292

,
   input                spc293_inst_done,
   input [63:0]         pc_w293

,
   input                spc294_inst_done,
   input [63:0]         pc_w294

,
   input                spc295_inst_done,
   input [63:0]         pc_w295

,
   input                spc296_inst_done,
   input [63:0]         pc_w296

,
   input                spc297_inst_done,
   input [63:0]         pc_w297

,
   input                spc298_inst_done,
   input [63:0]         pc_w298

,
   input                spc299_inst_done,
   input [63:0]         pc_w299

,
   input                spc300_inst_done,
   input [63:0]         pc_w300

,
   input                spc301_inst_done,
   input [63:0]         pc_w301

,
   input                spc302_inst_done,
   input [63:0]         pc_w302

,
   input                spc303_inst_done,
   input [63:0]         pc_w303

,
   input                spc304_inst_done,
   input [63:0]         pc_w304

,
   input                spc305_inst_done,
   input [63:0]         pc_w305

,
   input                spc306_inst_done,
   input [63:0]         pc_w306

,
   input                spc307_inst_done,
   input [63:0]         pc_w307

,
   input                spc308_inst_done,
   input [63:0]         pc_w308

,
   input                spc309_inst_done,
   input [63:0]         pc_w309

,
   input                spc310_inst_done,
   input [63:0]         pc_w310

,
   input                spc311_inst_done,
   input [63:0]         pc_w311

,
   input                spc312_inst_done,
   input [63:0]         pc_w312

,
   input                spc313_inst_done,
   input [63:0]         pc_w313

,
   input                spc314_inst_done,
   input [63:0]         pc_w314

,
   input                spc315_inst_done,
   input [63:0]         pc_w315

,
   input                spc316_inst_done,
   input [63:0]         pc_w316

,
   input                spc317_inst_done,
   input [63:0]         pc_w317

,
   input                spc318_inst_done,
   input [63:0]         pc_w318

,
   input                spc319_inst_done,
   input [63:0]         pc_w319

,
   input                spc320_inst_done,
   input [63:0]         pc_w320

,
   input                spc321_inst_done,
   input [63:0]         pc_w321

,
   input                spc322_inst_done,
   input [63:0]         pc_w322

,
   input                spc323_inst_done,
   input [63:0]         pc_w323

,
   input                spc324_inst_done,
   input [63:0]         pc_w324

,
   input                spc325_inst_done,
   input [63:0]         pc_w325

,
   input                spc326_inst_done,
   input [63:0]         pc_w326

,
   input                spc327_inst_done,
   input [63:0]         pc_w327

,
   input                spc328_inst_done,
   input [63:0]         pc_w328

,
   input                spc329_inst_done,
   input [63:0]         pc_w329

,
   input                spc330_inst_done,
   input [63:0]         pc_w330

,
   input                spc331_inst_done,
   input [63:0]         pc_w331

,
   input                spc332_inst_done,
   input [63:0]         pc_w332

,
   input                spc333_inst_done,
   input [63:0]         pc_w333

,
   input                spc334_inst_done,
   input [63:0]         pc_w334

,
   input                spc335_inst_done,
   input [63:0]         pc_w335

,
   input                spc336_inst_done,
   input [63:0]         pc_w336

,
   input                spc337_inst_done,
   input [63:0]         pc_w337

,
   input                spc338_inst_done,
   input [63:0]         pc_w338

,
   input                spc339_inst_done,
   input [63:0]         pc_w339

,
   input                spc340_inst_done,
   input [63:0]         pc_w340

,
   input                spc341_inst_done,
   input [63:0]         pc_w341

,
   input                spc342_inst_done,
   input [63:0]         pc_w342

,
   input                spc343_inst_done,
   input [63:0]         pc_w343

,
   input                spc344_inst_done,
   input [63:0]         pc_w344

,
   input                spc345_inst_done,
   input [63:0]         pc_w345

,
   input                spc346_inst_done,
   input [63:0]         pc_w346

,
   input                spc347_inst_done,
   input [63:0]         pc_w347

,
   input                spc348_inst_done,
   input [63:0]         pc_w348

,
   input                spc349_inst_done,
   input [63:0]         pc_w349

,
   input                spc350_inst_done,
   input [63:0]         pc_w350

,
   input                spc351_inst_done,
   input [63:0]         pc_w351

,
   input                spc352_inst_done,
   input [63:0]         pc_w352

,
   input                spc353_inst_done,
   input [63:0]         pc_w353

,
   input                spc354_inst_done,
   input [63:0]         pc_w354

,
   input                spc355_inst_done,
   input [63:0]         pc_w355

,
   input                spc356_inst_done,
   input [63:0]         pc_w356

,
   input                spc357_inst_done,
   input [63:0]         pc_w357

,
   input                spc358_inst_done,
   input [63:0]         pc_w358

,
   input                spc359_inst_done,
   input [63:0]         pc_w359

,
   input                spc360_inst_done,
   input [63:0]         pc_w360

,
   input                spc361_inst_done,
   input [63:0]         pc_w361

,
   input                spc362_inst_done,
   input [63:0]         pc_w362

,
   input                spc363_inst_done,
   input [63:0]         pc_w363

,
   input                spc364_inst_done,
   input [63:0]         pc_w364

,
   input                spc365_inst_done,
   input [63:0]         pc_w365

,
   input                spc366_inst_done,
   input [63:0]         pc_w366

,
   input                spc367_inst_done,
   input [63:0]         pc_w367

,
   input                spc368_inst_done,
   input [63:0]         pc_w368

,
   input                spc369_inst_done,
   input [63:0]         pc_w369

,
   input                spc370_inst_done,
   input [63:0]         pc_w370

,
   input                spc371_inst_done,
   input [63:0]         pc_w371

,
   input                spc372_inst_done,
   input [63:0]         pc_w372

,
   input                spc373_inst_done,
   input [63:0]         pc_w373

,
   input                spc374_inst_done,
   input [63:0]         pc_w374

,
   input                spc375_inst_done,
   input [63:0]         pc_w375

,
   input                spc376_inst_done,
   input [63:0]         pc_w376

,
   input                spc377_inst_done,
   input [63:0]         pc_w377

,
   input                spc378_inst_done,
   input [63:0]         pc_w378

,
   input                spc379_inst_done,
   input [63:0]         pc_w379

,
   input                spc380_inst_done,
   input [63:0]         pc_w380

,
   input                spc381_inst_done,
   input [63:0]         pc_w381

,
   input                spc382_inst_done,
   input [63:0]         pc_w382

,
   input                spc383_inst_done,
   input [63:0]         pc_w383

,
   input                spc384_inst_done,
   input [63:0]         pc_w384

,
   input                spc385_inst_done,
   input [63:0]         pc_w385

,
   input                spc386_inst_done,
   input [63:0]         pc_w386

,
   input                spc387_inst_done,
   input [63:0]         pc_w387

,
   input                spc388_inst_done,
   input [63:0]         pc_w388

,
   input                spc389_inst_done,
   input [63:0]         pc_w389

,
   input                spc390_inst_done,
   input [63:0]         pc_w390

,
   input                spc391_inst_done,
   input [63:0]         pc_w391

,
   input                spc392_inst_done,
   input [63:0]         pc_w392

,
   input                spc393_inst_done,
   input [63:0]         pc_w393

,
   input                spc394_inst_done,
   input [63:0]         pc_w394

,
   input                spc395_inst_done,
   input [63:0]         pc_w395

,
   input                spc396_inst_done,
   input [63:0]         pc_w396

,
   input                spc397_inst_done,
   input [63:0]         pc_w397

,
   input                spc398_inst_done,
   input [63:0]         pc_w398

,
   input                spc399_inst_done,
   input [63:0]         pc_w399

,
   input                spc400_inst_done,
   input [63:0]         pc_w400

,
   input                spc401_inst_done,
   input [63:0]         pc_w401

,
   input                spc402_inst_done,
   input [63:0]         pc_w402

,
   input                spc403_inst_done,
   input [63:0]         pc_w403

,
   input                spc404_inst_done,
   input [63:0]         pc_w404

,
   input                spc405_inst_done,
   input [63:0]         pc_w405

,
   input                spc406_inst_done,
   input [63:0]         pc_w406

,
   input                spc407_inst_done,
   input [63:0]         pc_w407

,
   input                spc408_inst_done,
   input [63:0]         pc_w408

,
   input                spc409_inst_done,
   input [63:0]         pc_w409

,
   input                spc410_inst_done,
   input [63:0]         pc_w410

,
   input                spc411_inst_done,
   input [63:0]         pc_w411

,
   input                spc412_inst_done,
   input [63:0]         pc_w412

,
   input                spc413_inst_done,
   input [63:0]         pc_w413

,
   input                spc414_inst_done,
   input [63:0]         pc_w414

,
   input                spc415_inst_done,
   input [63:0]         pc_w415

,
   input                spc416_inst_done,
   input [63:0]         pc_w416

,
   input                spc417_inst_done,
   input [63:0]         pc_w417

,
   input                spc418_inst_done,
   input [63:0]         pc_w418

,
   input                spc419_inst_done,
   input [63:0]         pc_w419

,
   input                spc420_inst_done,
   input [63:0]         pc_w420

,
   input                spc421_inst_done,
   input [63:0]         pc_w421

,
   input                spc422_inst_done,
   input [63:0]         pc_w422

,
   input                spc423_inst_done,
   input [63:0]         pc_w423

,
   input                spc424_inst_done,
   input [63:0]         pc_w424

,
   input                spc425_inst_done,
   input [63:0]         pc_w425

,
   input                spc426_inst_done,
   input [63:0]         pc_w426

,
   input                spc427_inst_done,
   input [63:0]         pc_w427

,
   input                spc428_inst_done,
   input [63:0]         pc_w428

,
   input                spc429_inst_done,
   input [63:0]         pc_w429

,
   input                spc430_inst_done,
   input [63:0]         pc_w430

,
   input                spc431_inst_done,
   input [63:0]         pc_w431

,
   input                spc432_inst_done,
   input [63:0]         pc_w432

,
   input                spc433_inst_done,
   input [63:0]         pc_w433

,
   input                spc434_inst_done,
   input [63:0]         pc_w434

,
   input                spc435_inst_done,
   input [63:0]         pc_w435

,
   input                spc436_inst_done,
   input [63:0]         pc_w436

,
   input                spc437_inst_done,
   input [63:0]         pc_w437

,
   input                spc438_inst_done,
   input [63:0]         pc_w438

,
   input                spc439_inst_done,
   input [63:0]         pc_w439

,
   input                spc440_inst_done,
   input [63:0]         pc_w440

,
   input                spc441_inst_done,
   input [63:0]         pc_w441

,
   input                spc442_inst_done,
   input [63:0]         pc_w442

,
   input                spc443_inst_done,
   input [63:0]         pc_w443

,
   input                spc444_inst_done,
   input [63:0]         pc_w444

,
   input                spc445_inst_done,
   input [63:0]         pc_w445

,
   input                spc446_inst_done,
   input [63:0]         pc_w446

,
   input                spc447_inst_done,
   input [63:0]         pc_w447

,
   input                spc448_inst_done,
   input [63:0]         pc_w448

,
   input                spc449_inst_done,
   input [63:0]         pc_w449

,
   input                spc450_inst_done,
   input [63:0]         pc_w450

,
   input                spc451_inst_done,
   input [63:0]         pc_w451

,
   input                spc452_inst_done,
   input [63:0]         pc_w452

,
   input                spc453_inst_done,
   input [63:0]         pc_w453

,
   input                spc454_inst_done,
   input [63:0]         pc_w454

,
   input                spc455_inst_done,
   input [63:0]         pc_w455

,
   input                spc456_inst_done,
   input [63:0]         pc_w456

,
   input                spc457_inst_done,
   input [63:0]         pc_w457

,
   input                spc458_inst_done,
   input [63:0]         pc_w458

,
   input                spc459_inst_done,
   input [63:0]         pc_w459

,
   input                spc460_inst_done,
   input [63:0]         pc_w460

,
   input                spc461_inst_done,
   input [63:0]         pc_w461

,
   input                spc462_inst_done,
   input [63:0]         pc_w462

,
   input                spc463_inst_done,
   input [63:0]         pc_w463

,
   input                spc464_inst_done,
   input [63:0]         pc_w464

,
   input                spc465_inst_done,
   input [63:0]         pc_w465

,
   input                spc466_inst_done,
   input [63:0]         pc_w466

,
   input                spc467_inst_done,
   input [63:0]         pc_w467

,
   input                spc468_inst_done,
   input [63:0]         pc_w468

,
   input                spc469_inst_done,
   input [63:0]         pc_w469

,
   input                spc470_inst_done,
   input [63:0]         pc_w470

,
   input                spc471_inst_done,
   input [63:0]         pc_w471

,
   input                spc472_inst_done,
   input [63:0]         pc_w472

,
   input                spc473_inst_done,
   input [63:0]         pc_w473

,
   input                spc474_inst_done,
   input [63:0]         pc_w474

,
   input                spc475_inst_done,
   input [63:0]         pc_w475

,
   input                spc476_inst_done,
   input [63:0]         pc_w476

,
   input                spc477_inst_done,
   input [63:0]         pc_w477

,
   input                spc478_inst_done,
   input [63:0]         pc_w478

,
   input                spc479_inst_done,
   input [63:0]         pc_w479

,
   input                spc480_inst_done,
   input [63:0]         pc_w480

,
   input                spc481_inst_done,
   input [63:0]         pc_w481

,
   input                spc482_inst_done,
   input [63:0]         pc_w482

,
   input                spc483_inst_done,
   input [63:0]         pc_w483

,
   input                spc484_inst_done,
   input [63:0]         pc_w484

,
   input                spc485_inst_done,
   input [63:0]         pc_w485

,
   input                spc486_inst_done,
   input [63:0]         pc_w486

,
   input                spc487_inst_done,
   input [63:0]         pc_w487

,
   input                spc488_inst_done,
   input [63:0]         pc_w488

,
   input                spc489_inst_done,
   input [63:0]         pc_w489

,
   input                spc490_inst_done,
   input [63:0]         pc_w490

,
   input                spc491_inst_done,
   input [63:0]         pc_w491

,
   input                spc492_inst_done,
   input [63:0]         pc_w492

,
   input                spc493_inst_done,
   input [63:0]         pc_w493

,
   input                spc494_inst_done,
   input [63:0]         pc_w494

,
   input                spc495_inst_done,
   input [63:0]         pc_w495

,
   input                spc496_inst_done,
   input [63:0]         pc_w496

,
   input                spc497_inst_done,
   input [63:0]         pc_w497

,
   input                spc498_inst_done,
   input [63:0]         pc_w498

,
   input                spc499_inst_done,
   input [63:0]         pc_w499

,
   input                spc500_inst_done,
   input [63:0]         pc_w500

,
   input                spc501_inst_done,
   input [63:0]         pc_w501

,
   input                spc502_inst_done,
   input [63:0]         pc_w502

,
   input                spc503_inst_done,
   input [63:0]         pc_w503

,
   input                spc504_inst_done,
   input [63:0]         pc_w504

,
   input                spc505_inst_done,
   input [63:0]         pc_w505

,
   input                spc506_inst_done,
   input [63:0]         pc_w506

,
   input                spc507_inst_done,
   input [63:0]         pc_w507

,
   input                spc508_inst_done,
   input [63:0]         pc_w508

,
   input                spc509_inst_done,
   input [63:0]         pc_w509

,
   input                spc510_inst_done,
   input [63:0]         pc_w510

,
   input                spc511_inst_done,
   input [63:0]         pc_w511

,
   input                spc512_inst_done,
   input [63:0]         pc_w512

,
   input                spc513_inst_done,
   input [63:0]         pc_w513

,
   input                spc514_inst_done,
   input [63:0]         pc_w514

,
   input                spc515_inst_done,
   input [63:0]         pc_w515

,
   input                spc516_inst_done,
   input [63:0]         pc_w516

,
   input                spc517_inst_done,
   input [63:0]         pc_w517

,
   input                spc518_inst_done,
   input [63:0]         pc_w518

,
   input                spc519_inst_done,
   input [63:0]         pc_w519

,
   input                spc520_inst_done,
   input [63:0]         pc_w520

,
   input                spc521_inst_done,
   input [63:0]         pc_w521

,
   input                spc522_inst_done,
   input [63:0]         pc_w522

,
   input                spc523_inst_done,
   input [63:0]         pc_w523

,
   input                spc524_inst_done,
   input [63:0]         pc_w524

,
   input                spc525_inst_done,
   input [63:0]         pc_w525

,
   input                spc526_inst_done,
   input [63:0]         pc_w526

,
   input                spc527_inst_done,
   input [63:0]         pc_w527

,
   input                spc528_inst_done,
   input [63:0]         pc_w528

,
   input                spc529_inst_done,
   input [63:0]         pc_w529

,
   input                spc530_inst_done,
   input [63:0]         pc_w530

,
   input                spc531_inst_done,
   input [63:0]         pc_w531

,
   input                spc532_inst_done,
   input [63:0]         pc_w532

,
   input                spc533_inst_done,
   input [63:0]         pc_w533

,
   input                spc534_inst_done,
   input [63:0]         pc_w534

,
   input                spc535_inst_done,
   input [63:0]         pc_w535

,
   input                spc536_inst_done,
   input [63:0]         pc_w536

,
   input                spc537_inst_done,
   input [63:0]         pc_w537

,
   input                spc538_inst_done,
   input [63:0]         pc_w538

,
   input                spc539_inst_done,
   input [63:0]         pc_w539

,
   input                spc540_inst_done,
   input [63:0]         pc_w540

,
   input                spc541_inst_done,
   input [63:0]         pc_w541

,
   input                spc542_inst_done,
   input [63:0]         pc_w542

,
   input                spc543_inst_done,
   input [63:0]         pc_w543

,
   input                spc544_inst_done,
   input [63:0]         pc_w544

,
   input                spc545_inst_done,
   input [63:0]         pc_w545

,
   input                spc546_inst_done,
   input [63:0]         pc_w546

,
   input                spc547_inst_done,
   input [63:0]         pc_w547

,
   input                spc548_inst_done,
   input [63:0]         pc_w548

,
   input                spc549_inst_done,
   input [63:0]         pc_w549

,
   input                spc550_inst_done,
   input [63:0]         pc_w550

,
   input                spc551_inst_done,
   input [63:0]         pc_w551

,
   input                spc552_inst_done,
   input [63:0]         pc_w552

,
   input                spc553_inst_done,
   input [63:0]         pc_w553

,
   input                spc554_inst_done,
   input [63:0]         pc_w554

,
   input                spc555_inst_done,
   input [63:0]         pc_w555

,
   input                spc556_inst_done,
   input [63:0]         pc_w556

,
   input                spc557_inst_done,
   input [63:0]         pc_w557

,
   input                spc558_inst_done,
   input [63:0]         pc_w558

,
   input                spc559_inst_done,
   input [63:0]         pc_w559

,
   input                spc560_inst_done,
   input [63:0]         pc_w560

,
   input                spc561_inst_done,
   input [63:0]         pc_w561

,
   input                spc562_inst_done,
   input [63:0]         pc_w562

,
   input                spc563_inst_done,
   input [63:0]         pc_w563

,
   input                spc564_inst_done,
   input [63:0]         pc_w564

,
   input                spc565_inst_done,
   input [63:0]         pc_w565

,
   input                spc566_inst_done,
   input [63:0]         pc_w566

,
   input                spc567_inst_done,
   input [63:0]         pc_w567

,
   input                spc568_inst_done,
   input [63:0]         pc_w568

,
   input                spc569_inst_done,
   input [63:0]         pc_w569

,
   input                spc570_inst_done,
   input [63:0]         pc_w570

,
   input                spc571_inst_done,
   input [63:0]         pc_w571

,
   input                spc572_inst_done,
   input [63:0]         pc_w572

,
   input                spc573_inst_done,
   input [63:0]         pc_w573

,
   input                spc574_inst_done,
   input [63:0]         pc_w574

,
   input                spc575_inst_done,
   input [63:0]         pc_w575

,
   input                spc576_inst_done,
   input [63:0]         pc_w576

,
   input                spc577_inst_done,
   input [63:0]         pc_w577

,
   input                spc578_inst_done,
   input [63:0]         pc_w578

,
   input                spc579_inst_done,
   input [63:0]         pc_w579

,
   input                spc580_inst_done,
   input [63:0]         pc_w580

,
   input                spc581_inst_done,
   input [63:0]         pc_w581

,
   input                spc582_inst_done,
   input [63:0]         pc_w582

,
   input                spc583_inst_done,
   input [63:0]         pc_w583

,
   input                spc584_inst_done,
   input [63:0]         pc_w584

,
   input                spc585_inst_done,
   input [63:0]         pc_w585

,
   input                spc586_inst_done,
   input [63:0]         pc_w586

,
   input                spc587_inst_done,
   input [63:0]         pc_w587

,
   input                spc588_inst_done,
   input [63:0]         pc_w588

,
   input                spc589_inst_done,
   input [63:0]         pc_w589

,
   input                spc590_inst_done,
   input [63:0]         pc_w590

,
   input                spc591_inst_done,
   input [63:0]         pc_w591

,
   input                spc592_inst_done,
   input [63:0]         pc_w592

,
   input                spc593_inst_done,
   input [63:0]         pc_w593

,
   input                spc594_inst_done,
   input [63:0]         pc_w594

,
   input                spc595_inst_done,
   input [63:0]         pc_w595

,
   input                spc596_inst_done,
   input [63:0]         pc_w596

,
   input                spc597_inst_done,
   input [63:0]         pc_w597

,
   input                spc598_inst_done,
   input [63:0]         pc_w598

,
   input                spc599_inst_done,
   input [63:0]         pc_w599

,
   input                spc600_inst_done,
   input [63:0]         pc_w600

,
   input                spc601_inst_done,
   input [63:0]         pc_w601

,
   input                spc602_inst_done,
   input [63:0]         pc_w602

,
   input                spc603_inst_done,
   input [63:0]         pc_w603

,
   input                spc604_inst_done,
   input [63:0]         pc_w604

,
   input                spc605_inst_done,
   input [63:0]         pc_w605

,
   input                spc606_inst_done,
   input [63:0]         pc_w606

,
   input                spc607_inst_done,
   input [63:0]         pc_w607

,
   input                spc608_inst_done,
   input [63:0]         pc_w608

,
   input                spc609_inst_done,
   input [63:0]         pc_w609

,
   input                spc610_inst_done,
   input [63:0]         pc_w610

,
   input                spc611_inst_done,
   input [63:0]         pc_w611

,
   input                spc612_inst_done,
   input [63:0]         pc_w612

,
   input                spc613_inst_done,
   input [63:0]         pc_w613

,
   input                spc614_inst_done,
   input [63:0]         pc_w614

,
   input                spc615_inst_done,
   input [63:0]         pc_w615

,
   input                spc616_inst_done,
   input [63:0]         pc_w616

,
   input                spc617_inst_done,
   input [63:0]         pc_w617

,
   input                spc618_inst_done,
   input [63:0]         pc_w618

,
   input                spc619_inst_done,
   input [63:0]         pc_w619

,
   input                spc620_inst_done,
   input [63:0]         pc_w620

,
   input                spc621_inst_done,
   input [63:0]         pc_w621

,
   input                spc622_inst_done,
   input [63:0]         pc_w622

,
   input                spc623_inst_done,
   input [63:0]         pc_w623

,
   input                spc624_inst_done,
   input [63:0]         pc_w624

,
   input                spc625_inst_done,
   input [63:0]         pc_w625

,
   input                spc626_inst_done,
   input [63:0]         pc_w626

,
   input                spc627_inst_done,
   input [63:0]         pc_w627

,
   input                spc628_inst_done,
   input [63:0]         pc_w628

,
   input                spc629_inst_done,
   input [63:0]         pc_w629

,
   input                spc630_inst_done,
   input [63:0]         pc_w630

,
   input                spc631_inst_done,
   input [63:0]         pc_w631

,
   input                spc632_inst_done,
   input [63:0]         pc_w632

,
   input                spc633_inst_done,
   input [63:0]         pc_w633

,
   input                spc634_inst_done,
   input [63:0]         pc_w634

,
   input                spc635_inst_done,
   input [63:0]         pc_w635

,
   input                spc636_inst_done,
   input [63:0]         pc_w636

,
   input                spc637_inst_done,
   input [63:0]         pc_w637

,
   input                spc638_inst_done,
   input [63:0]         pc_w638

,
   input                spc639_inst_done,
   input [63:0]         pc_w639

,
   input                spc640_inst_done,
   input [63:0]         pc_w640

,
   input                spc641_inst_done,
   input [63:0]         pc_w641

,
   input                spc642_inst_done,
   input [63:0]         pc_w642

,
   input                spc643_inst_done,
   input [63:0]         pc_w643

,
   input                spc644_inst_done,
   input [63:0]         pc_w644

,
   input                spc645_inst_done,
   input [63:0]         pc_w645

,
   input                spc646_inst_done,
   input [63:0]         pc_w646

,
   input                spc647_inst_done,
   input [63:0]         pc_w647

,
   input                spc648_inst_done,
   input [63:0]         pc_w648

,
   input                spc649_inst_done,
   input [63:0]         pc_w649

,
   input                spc650_inst_done,
   input [63:0]         pc_w650

,
   input                spc651_inst_done,
   input [63:0]         pc_w651

,
   input                spc652_inst_done,
   input [63:0]         pc_w652

,
   input                spc653_inst_done,
   input [63:0]         pc_w653

,
   input                spc654_inst_done,
   input [63:0]         pc_w654

,
   input                spc655_inst_done,
   input [63:0]         pc_w655

,
   input                spc656_inst_done,
   input [63:0]         pc_w656

,
   input                spc657_inst_done,
   input [63:0]         pc_w657

,
   input                spc658_inst_done,
   input [63:0]         pc_w658

,
   input                spc659_inst_done,
   input [63:0]         pc_w659

,
   input                spc660_inst_done,
   input [63:0]         pc_w660

,
   input                spc661_inst_done,
   input [63:0]         pc_w661

,
   input                spc662_inst_done,
   input [63:0]         pc_w662

,
   input                spc663_inst_done,
   input [63:0]         pc_w663

,
   input                spc664_inst_done,
   input [63:0]         pc_w664

,
   input                spc665_inst_done,
   input [63:0]         pc_w665

,
   input                spc666_inst_done,
   input [63:0]         pc_w666

,
   input                spc667_inst_done,
   input [63:0]         pc_w667

,
   input                spc668_inst_done,
   input [63:0]         pc_w668

,
   input                spc669_inst_done,
   input [63:0]         pc_w669

,
   input                spc670_inst_done,
   input [63:0]         pc_w670

,
   input                spc671_inst_done,
   input [63:0]         pc_w671

,
   input                spc672_inst_done,
   input [63:0]         pc_w672

,
   input                spc673_inst_done,
   input [63:0]         pc_w673

,
   input                spc674_inst_done,
   input [63:0]         pc_w674

,
   input                spc675_inst_done,
   input [63:0]         pc_w675

,
   input                spc676_inst_done,
   input [63:0]         pc_w676

,
   input                spc677_inst_done,
   input [63:0]         pc_w677

,
   input                spc678_inst_done,
   input [63:0]         pc_w678

,
   input                spc679_inst_done,
   input [63:0]         pc_w679

,
   input                spc680_inst_done,
   input [63:0]         pc_w680

,
   input                spc681_inst_done,
   input [63:0]         pc_w681

,
   input                spc682_inst_done,
   input [63:0]         pc_w682

,
   input                spc683_inst_done,
   input [63:0]         pc_w683

,
   input                spc684_inst_done,
   input [63:0]         pc_w684

,
   input                spc685_inst_done,
   input [63:0]         pc_w685

,
   input                spc686_inst_done,
   input [63:0]         pc_w686

,
   input                spc687_inst_done,
   input [63:0]         pc_w687

,
   input                spc688_inst_done,
   input [63:0]         pc_w688

,
   input                spc689_inst_done,
   input [63:0]         pc_w689

,
   input                spc690_inst_done,
   input [63:0]         pc_w690

,
   input                spc691_inst_done,
   input [63:0]         pc_w691

,
   input                spc692_inst_done,
   input [63:0]         pc_w692

,
   input                spc693_inst_done,
   input [63:0]         pc_w693

,
   input                spc694_inst_done,
   input [63:0]         pc_w694

,
   input                spc695_inst_done,
   input [63:0]         pc_w695

,
   input                spc696_inst_done,
   input [63:0]         pc_w696

,
   input                spc697_inst_done,
   input [63:0]         pc_w697

,
   input                spc698_inst_done,
   input [63:0]         pc_w698

,
   input                spc699_inst_done,
   input [63:0]         pc_w699

,
   input                spc700_inst_done,
   input [63:0]         pc_w700

,
   input                spc701_inst_done,
   input [63:0]         pc_w701

,
   input                spc702_inst_done,
   input [63:0]         pc_w702

,
   input                spc703_inst_done,
   input [63:0]         pc_w703

,
   input                spc704_inst_done,
   input [63:0]         pc_w704

,
   input                spc705_inst_done,
   input [63:0]         pc_w705

,
   input                spc706_inst_done,
   input [63:0]         pc_w706

,
   input                spc707_inst_done,
   input [63:0]         pc_w707

,
   input                spc708_inst_done,
   input [63:0]         pc_w708

,
   input                spc709_inst_done,
   input [63:0]         pc_w709

,
   input                spc710_inst_done,
   input [63:0]         pc_w710

,
   input                spc711_inst_done,
   input [63:0]         pc_w711

,
   input                spc712_inst_done,
   input [63:0]         pc_w712

,
   input                spc713_inst_done,
   input [63:0]         pc_w713

,
   input                spc714_inst_done,
   input [63:0]         pc_w714

,
   input                spc715_inst_done,
   input [63:0]         pc_w715

,
   input                spc716_inst_done,
   input [63:0]         pc_w716

,
   input                spc717_inst_done,
   input [63:0]         pc_w717

,
   input                spc718_inst_done,
   input [63:0]         pc_w718

,
   input                spc719_inst_done,
   input [63:0]         pc_w719

,
   input                spc720_inst_done,
   input [63:0]         pc_w720

,
   input                spc721_inst_done,
   input [63:0]         pc_w721

,
   input                spc722_inst_done,
   input [63:0]         pc_w722

,
   input                spc723_inst_done,
   input [63:0]         pc_w723

,
   input                spc724_inst_done,
   input [63:0]         pc_w724

,
   input                spc725_inst_done,
   input [63:0]         pc_w725

,
   input                spc726_inst_done,
   input [63:0]         pc_w726

,
   input                spc727_inst_done,
   input [63:0]         pc_w727

,
   input                spc728_inst_done,
   input [63:0]         pc_w728

,
   input                spc729_inst_done,
   input [63:0]         pc_w729

,
   input                spc730_inst_done,
   input [63:0]         pc_w730

,
   input                spc731_inst_done,
   input [63:0]         pc_w731

,
   input                spc732_inst_done,
   input [63:0]         pc_w732

,
   input                spc733_inst_done,
   input [63:0]         pc_w733

,
   input                spc734_inst_done,
   input [63:0]         pc_w734

,
   input                spc735_inst_done,
   input [63:0]         pc_w735

,
   input                spc736_inst_done,
   input [63:0]         pc_w736

,
   input                spc737_inst_done,
   input [63:0]         pc_w737

,
   input                spc738_inst_done,
   input [63:0]         pc_w738

,
   input                spc739_inst_done,
   input [63:0]         pc_w739

,
   input                spc740_inst_done,
   input [63:0]         pc_w740

,
   input                spc741_inst_done,
   input [63:0]         pc_w741

,
   input                spc742_inst_done,
   input [63:0]         pc_w742

,
   input                spc743_inst_done,
   input [63:0]         pc_w743

,
   input                spc744_inst_done,
   input [63:0]         pc_w744

,
   input                spc745_inst_done,
   input [63:0]         pc_w745

,
   input                spc746_inst_done,
   input [63:0]         pc_w746

,
   input                spc747_inst_done,
   input [63:0]         pc_w747

,
   input                spc748_inst_done,
   input [63:0]         pc_w748

,
   input                spc749_inst_done,
   input [63:0]         pc_w749

,
   input                spc750_inst_done,
   input [63:0]         pc_w750

,
   input                spc751_inst_done,
   input [63:0]         pc_w751

,
   input                spc752_inst_done,
   input [63:0]         pc_w752

,
   input                spc753_inst_done,
   input [63:0]         pc_w753

,
   input                spc754_inst_done,
   input [63:0]         pc_w754

,
   input                spc755_inst_done,
   input [63:0]         pc_w755

,
   input                spc756_inst_done,
   input [63:0]         pc_w756

,
   input                spc757_inst_done,
   input [63:0]         pc_w757

,
   input                spc758_inst_done,
   input [63:0]         pc_w758

,
   input                spc759_inst_done,
   input [63:0]         pc_w759

,
   input                spc760_inst_done,
   input [63:0]         pc_w760

,
   input                spc761_inst_done,
   input [63:0]         pc_w761

,
   input                spc762_inst_done,
   input [63:0]         pc_w762

,
   input                spc763_inst_done,
   input [63:0]         pc_w763

,
   input                spc764_inst_done,
   input [63:0]         pc_w764

,
   input                spc765_inst_done,
   input [63:0]         pc_w765

,
   input                spc766_inst_done,
   input [63:0]         pc_w766

,
   input                spc767_inst_done,
   input [63:0]         pc_w767

,
   input                spc768_inst_done,
   input [63:0]         pc_w768

,
   input                spc769_inst_done,
   input [63:0]         pc_w769

,
   input                spc770_inst_done,
   input [63:0]         pc_w770

,
   input                spc771_inst_done,
   input [63:0]         pc_w771

,
   input                spc772_inst_done,
   input [63:0]         pc_w772

,
   input                spc773_inst_done,
   input [63:0]         pc_w773

,
   input                spc774_inst_done,
   input [63:0]         pc_w774

,
   input                spc775_inst_done,
   input [63:0]         pc_w775

,
   input                spc776_inst_done,
   input [63:0]         pc_w776

,
   input                spc777_inst_done,
   input [63:0]         pc_w777

,
   input                spc778_inst_done,
   input [63:0]         pc_w778

,
   input                spc779_inst_done,
   input [63:0]         pc_w779

,
   input                spc780_inst_done,
   input [63:0]         pc_w780

,
   input                spc781_inst_done,
   input [63:0]         pc_w781

,
   input                spc782_inst_done,
   input [63:0]         pc_w782

,
   input                spc783_inst_done,
   input [63:0]         pc_w783

,
   input                spc784_inst_done,
   input [63:0]         pc_w784

,
   input                spc785_inst_done,
   input [63:0]         pc_w785

,
   input                spc786_inst_done,
   input [63:0]         pc_w786

,
   input                spc787_inst_done,
   input [63:0]         pc_w787

,
   input                spc788_inst_done,
   input [63:0]         pc_w788

,
   input                spc789_inst_done,
   input [63:0]         pc_w789

,
   input                spc790_inst_done,
   input [63:0]         pc_w790

,
   input                spc791_inst_done,
   input [63:0]         pc_w791

,
   input                spc792_inst_done,
   input [63:0]         pc_w792

,
   input                spc793_inst_done,
   input [63:0]         pc_w793

,
   input                spc794_inst_done,
   input [63:0]         pc_w794

,
   input                spc795_inst_done,
   input [63:0]         pc_w795

,
   input                spc796_inst_done,
   input [63:0]         pc_w796

,
   input                spc797_inst_done,
   input [63:0]         pc_w797

,
   input                spc798_inst_done,
   input [63:0]         pc_w798

,
   input                spc799_inst_done,
   input [63:0]         pc_w799

,
   input                spc800_inst_done,
   input [63:0]         pc_w800

,
   input                spc801_inst_done,
   input [63:0]         pc_w801

,
   input                spc802_inst_done,
   input [63:0]         pc_w802

,
   input                spc803_inst_done,
   input [63:0]         pc_w803

,
   input                spc804_inst_done,
   input [63:0]         pc_w804

,
   input                spc805_inst_done,
   input [63:0]         pc_w805

,
   input                spc806_inst_done,
   input [63:0]         pc_w806

,
   input                spc807_inst_done,
   input [63:0]         pc_w807

,
   input                spc808_inst_done,
   input [63:0]         pc_w808

,
   input                spc809_inst_done,
   input [63:0]         pc_w809

,
   input                spc810_inst_done,
   input [63:0]         pc_w810

,
   input                spc811_inst_done,
   input [63:0]         pc_w811

,
   input                spc812_inst_done,
   input [63:0]         pc_w812

,
   input                spc813_inst_done,
   input [63:0]         pc_w813

,
   input                spc814_inst_done,
   input [63:0]         pc_w814

,
   input                spc815_inst_done,
   input [63:0]         pc_w815

,
   input                spc816_inst_done,
   input [63:0]         pc_w816

,
   input                spc817_inst_done,
   input [63:0]         pc_w817

,
   input                spc818_inst_done,
   input [63:0]         pc_w818

,
   input                spc819_inst_done,
   input [63:0]         pc_w819

,
   input                spc820_inst_done,
   input [63:0]         pc_w820

,
   input                spc821_inst_done,
   input [63:0]         pc_w821

,
   input                spc822_inst_done,
   input [63:0]         pc_w822

,
   input                spc823_inst_done,
   input [63:0]         pc_w823

,
   input                spc824_inst_done,
   input [63:0]         pc_w824

,
   input                spc825_inst_done,
   input [63:0]         pc_w825

,
   input                spc826_inst_done,
   input [63:0]         pc_w826

,
   input                spc827_inst_done,
   input [63:0]         pc_w827

,
   input                spc828_inst_done,
   input [63:0]         pc_w828

,
   input                spc829_inst_done,
   input [63:0]         pc_w829

,
   input                spc830_inst_done,
   input [63:0]         pc_w830

,
   input                spc831_inst_done,
   input [63:0]         pc_w831

,
   input                spc832_inst_done,
   input [63:0]         pc_w832

,
   input                spc833_inst_done,
   input [63:0]         pc_w833

,
   input                spc834_inst_done,
   input [63:0]         pc_w834

,
   input                spc835_inst_done,
   input [63:0]         pc_w835

,
   input                spc836_inst_done,
   input [63:0]         pc_w836

,
   input                spc837_inst_done,
   input [63:0]         pc_w837

,
   input                spc838_inst_done,
   input [63:0]         pc_w838

,
   input                spc839_inst_done,
   input [63:0]         pc_w839

,
   input                spc840_inst_done,
   input [63:0]         pc_w840

,
   input                spc841_inst_done,
   input [63:0]         pc_w841

,
   input                spc842_inst_done,
   input [63:0]         pc_w842

,
   input                spc843_inst_done,
   input [63:0]         pc_w843

,
   input                spc844_inst_done,
   input [63:0]         pc_w844

,
   input                spc845_inst_done,
   input [63:0]         pc_w845

,
   input                spc846_inst_done,
   input [63:0]         pc_w846

,
   input                spc847_inst_done,
   input [63:0]         pc_w847

,
   input                spc848_inst_done,
   input [63:0]         pc_w848

,
   input                spc849_inst_done,
   input [63:0]         pc_w849

,
   input                spc850_inst_done,
   input [63:0]         pc_w850

,
   input                spc851_inst_done,
   input [63:0]         pc_w851

,
   input                spc852_inst_done,
   input [63:0]         pc_w852

,
   input                spc853_inst_done,
   input [63:0]         pc_w853

,
   input                spc854_inst_done,
   input [63:0]         pc_w854

,
   input                spc855_inst_done,
   input [63:0]         pc_w855

,
   input                spc856_inst_done,
   input [63:0]         pc_w856

,
   input                spc857_inst_done,
   input [63:0]         pc_w857

,
   input                spc858_inst_done,
   input [63:0]         pc_w858

,
   input                spc859_inst_done,
   input [63:0]         pc_w859

,
   input                spc860_inst_done,
   input [63:0]         pc_w860

,
   input                spc861_inst_done,
   input [63:0]         pc_w861

,
   input                spc862_inst_done,
   input [63:0]         pc_w862

,
   input                spc863_inst_done,
   input [63:0]         pc_w863

,
   input                spc864_inst_done,
   input [63:0]         pc_w864

,
   input                spc865_inst_done,
   input [63:0]         pc_w865

,
   input                spc866_inst_done,
   input [63:0]         pc_w866

,
   input                spc867_inst_done,
   input [63:0]         pc_w867

,
   input                spc868_inst_done,
   input [63:0]         pc_w868

,
   input                spc869_inst_done,
   input [63:0]         pc_w869

,
   input                spc870_inst_done,
   input [63:0]         pc_w870

,
   input                spc871_inst_done,
   input [63:0]         pc_w871

,
   input                spc872_inst_done,
   input [63:0]         pc_w872

,
   input                spc873_inst_done,
   input [63:0]         pc_w873

,
   input                spc874_inst_done,
   input [63:0]         pc_w874

,
   input                spc875_inst_done,
   input [63:0]         pc_w875

,
   input                spc876_inst_done,
   input [63:0]         pc_w876

,
   input                spc877_inst_done,
   input [63:0]         pc_w877

,
   input                spc878_inst_done,
   input [63:0]         pc_w878

,
   input                spc879_inst_done,
   input [63:0]         pc_w879

,
   input                spc880_inst_done,
   input [63:0]         pc_w880

,
   input                spc881_inst_done,
   input [63:0]         pc_w881

,
   input                spc882_inst_done,
   input [63:0]         pc_w882

,
   input                spc883_inst_done,
   input [63:0]         pc_w883

,
   input                spc884_inst_done,
   input [63:0]         pc_w884

,
   input                spc885_inst_done,
   input [63:0]         pc_w885

,
   input                spc886_inst_done,
   input [63:0]         pc_w886

,
   input                spc887_inst_done,
   input [63:0]         pc_w887

,
   input                spc888_inst_done,
   input [63:0]         pc_w888

,
   input                spc889_inst_done,
   input [63:0]         pc_w889

,
   input                spc890_inst_done,
   input [63:0]         pc_w890

,
   input                spc891_inst_done,
   input [63:0]         pc_w891

,
   input                spc892_inst_done,
   input [63:0]         pc_w892

,
   input                spc893_inst_done,
   input [63:0]         pc_w893

,
   input                spc894_inst_done,
   input [63:0]         pc_w894

,
   input                spc895_inst_done,
   input [63:0]         pc_w895

,
   input                spc896_inst_done,
   input [63:0]         pc_w896

,
   input                spc897_inst_done,
   input [63:0]         pc_w897

,
   input                spc898_inst_done,
   input [63:0]         pc_w898

,
   input                spc899_inst_done,
   input [63:0]         pc_w899

,
   input                spc900_inst_done,
   input [63:0]         pc_w900

,
   input                spc901_inst_done,
   input [63:0]         pc_w901

,
   input                spc902_inst_done,
   input [63:0]         pc_w902

,
   input                spc903_inst_done,
   input [63:0]         pc_w903

,
   input                spc904_inst_done,
   input [63:0]         pc_w904

,
   input                spc905_inst_done,
   input [63:0]         pc_w905

,
   input                spc906_inst_done,
   input [63:0]         pc_w906

,
   input                spc907_inst_done,
   input [63:0]         pc_w907

,
   input                spc908_inst_done,
   input [63:0]         pc_w908

,
   input                spc909_inst_done,
   input [63:0]         pc_w909

,
   input                spc910_inst_done,
   input [63:0]         pc_w910

,
   input                spc911_inst_done,
   input [63:0]         pc_w911

,
   input                spc912_inst_done,
   input [63:0]         pc_w912

,
   input                spc913_inst_done,
   input [63:0]         pc_w913

,
   input                spc914_inst_done,
   input [63:0]         pc_w914

,
   input                spc915_inst_done,
   input [63:0]         pc_w915

,
   input                spc916_inst_done,
   input [63:0]         pc_w916

,
   input                spc917_inst_done,
   input [63:0]         pc_w917

,
   input                spc918_inst_done,
   input [63:0]         pc_w918

,
   input                spc919_inst_done,
   input [63:0]         pc_w919

,
   input                spc920_inst_done,
   input [63:0]         pc_w920

,
   input                spc921_inst_done,
   input [63:0]         pc_w921

,
   input                spc922_inst_done,
   input [63:0]         pc_w922

,
   input                spc923_inst_done,
   input [63:0]         pc_w923

,
   input                spc924_inst_done,
   input [63:0]         pc_w924

,
   input                spc925_inst_done,
   input [63:0]         pc_w925

,
   input                spc926_inst_done,
   input [63:0]         pc_w926

,
   input                spc927_inst_done,
   input [63:0]         pc_w927

,
   input                spc928_inst_done,
   input [63:0]         pc_w928

,
   input                spc929_inst_done,
   input [63:0]         pc_w929

,
   input                spc930_inst_done,
   input [63:0]         pc_w930

,
   input                spc931_inst_done,
   input [63:0]         pc_w931

,
   input                spc932_inst_done,
   input [63:0]         pc_w932

,
   input                spc933_inst_done,
   input [63:0]         pc_w933

,
   input                spc934_inst_done,
   input [63:0]         pc_w934

,
   input                spc935_inst_done,
   input [63:0]         pc_w935

,
   input                spc936_inst_done,
   input [63:0]         pc_w936

,
   input                spc937_inst_done,
   input [63:0]         pc_w937

,
   input                spc938_inst_done,
   input [63:0]         pc_w938

,
   input                spc939_inst_done,
   input [63:0]         pc_w939

,
   input                spc940_inst_done,
   input [63:0]         pc_w940

,
   input                spc941_inst_done,
   input [63:0]         pc_w941

,
   input                spc942_inst_done,
   input [63:0]         pc_w942

,
   input                spc943_inst_done,
   input [63:0]         pc_w943

,
   input                spc944_inst_done,
   input [63:0]         pc_w944

,
   input                spc945_inst_done,
   input [63:0]         pc_w945

,
   input                spc946_inst_done,
   input [63:0]         pc_w946

,
   input                spc947_inst_done,
   input [63:0]         pc_w947

,
   input                spc948_inst_done,
   input [63:0]         pc_w948

,
   input                spc949_inst_done,
   input [63:0]         pc_w949

,
   input                spc950_inst_done,
   input [63:0]         pc_w950

,
   input                spc951_inst_done,
   input [63:0]         pc_w951

,
   input                spc952_inst_done,
   input [63:0]         pc_w952

,
   input                spc953_inst_done,
   input [63:0]         pc_w953

,
   input                spc954_inst_done,
   input [63:0]         pc_w954

,
   input                spc955_inst_done,
   input [63:0]         pc_w955

,
   input                spc956_inst_done,
   input [63:0]         pc_w956

,
   input                spc957_inst_done,
   input [63:0]         pc_w957

,
   input                spc958_inst_done,
   input [63:0]         pc_w958

,
   input                spc959_inst_done,
   input [63:0]         pc_w959

,
   input                spc960_inst_done,
   input [63:0]         pc_w960

,
   input                spc961_inst_done,
   input [63:0]         pc_w961

,
   input                spc962_inst_done,
   input [63:0]         pc_w962

,
   input                spc963_inst_done,
   input [63:0]         pc_w963

,
   input                spc964_inst_done,
   input [63:0]         pc_w964

,
   input                spc965_inst_done,
   input [63:0]         pc_w965

,
   input                spc966_inst_done,
   input [63:0]         pc_w966

,
   input                spc967_inst_done,
   input [63:0]         pc_w967

,
   input                spc968_inst_done,
   input [63:0]         pc_w968

,
   input                spc969_inst_done,
   input [63:0]         pc_w969

,
   input                spc970_inst_done,
   input [63:0]         pc_w970

,
   input                spc971_inst_done,
   input [63:0]         pc_w971

,
   input                spc972_inst_done,
   input [63:0]         pc_w972

,
   input                spc973_inst_done,
   input [63:0]         pc_w973

,
   input                spc974_inst_done,
   input [63:0]         pc_w974

,
   input                spc975_inst_done,
   input [63:0]         pc_w975

,
   input                spc976_inst_done,
   input [63:0]         pc_w976

,
   input                spc977_inst_done,
   input [63:0]         pc_w977

,
   input                spc978_inst_done,
   input [63:0]         pc_w978

,
   input                spc979_inst_done,
   input [63:0]         pc_w979

,
   input                spc980_inst_done,
   input [63:0]         pc_w980

,
   input                spc981_inst_done,
   input [63:0]         pc_w981

,
   input                spc982_inst_done,
   input [63:0]         pc_w982

,
   input                spc983_inst_done,
   input [63:0]         pc_w983

,
   input                spc984_inst_done,
   input [63:0]         pc_w984

,
   input                spc985_inst_done,
   input [63:0]         pc_w985

,
   input                spc986_inst_done,
   input [63:0]         pc_w986

,
   input                spc987_inst_done,
   input [63:0]         pc_w987

,
   input                spc988_inst_done,
   input [63:0]         pc_w988

,
   input                spc989_inst_done,
   input [63:0]         pc_w989

,
   input                spc990_inst_done,
   input [63:0]         pc_w990

,
   input                spc991_inst_done,
   input [63:0]         pc_w991

,
   input                spc992_inst_done,
   input [63:0]         pc_w992

,
   input                spc993_inst_done,
   input [63:0]         pc_w993

,
   input                spc994_inst_done,
   input [63:0]         pc_w994

,
   input                spc995_inst_done,
   input [63:0]         pc_w995

,
   input                spc996_inst_done,
   input [63:0]         pc_w996

,
   input                spc997_inst_done,
   input [63:0]         pc_w997

,
   input                spc998_inst_done,
   input [63:0]         pc_w998

,
   input                spc999_inst_done,
   input [63:0]         pc_w999

,
   input                spc1000_inst_done,
   input [63:0]         pc_w1000

,
   input                spc1001_inst_done,
   input [63:0]         pc_w1001

,
   input                spc1002_inst_done,
   input [63:0]         pc_w1002

,
   input                spc1003_inst_done,
   input [63:0]         pc_w1003

,
   input                spc1004_inst_done,
   input [63:0]         pc_w1004

,
   input                spc1005_inst_done,
   input [63:0]         pc_w1005

,
   input                spc1006_inst_done,
   input [63:0]         pc_w1006

,
   input                spc1007_inst_done,
   input [63:0]         pc_w1007

,
   input                spc1008_inst_done,
   input [63:0]         pc_w1008

,
   input                spc1009_inst_done,
   input [63:0]         pc_w1009

,
   input                spc1010_inst_done,
   input [63:0]         pc_w1010

,
   input                spc1011_inst_done,
   input [63:0]         pc_w1011

,
   input                spc1012_inst_done,
   input [63:0]         pc_w1012

,
   input                spc1013_inst_done,
   input [63:0]         pc_w1013

,
   input                spc1014_inst_done,
   input [63:0]         pc_w1014

,
   input                spc1015_inst_done,
   input [63:0]         pc_w1015

,
   input                spc1016_inst_done,
   input [63:0]         pc_w1016

,
   input                spc1017_inst_done,
   input [63:0]         pc_w1017

,
   input                spc1018_inst_done,
   input [63:0]         pc_w1018

,
   input                spc1019_inst_done,
   input [63:0]         pc_w1019

,
   input                spc1020_inst_done,
   input [63:0]         pc_w1020

,
   input                spc1021_inst_done,
   input [63:0]         pc_w1021

,
   input                spc1022_inst_done,
   input [63:0]         pc_w1022

,
   input                spc1023_inst_done,
   input [63:0]         pc_w1023



);
//temp. memory.
reg [`CPX_WIDTH-1:0] 	    fake_iob_out_data;

wire [`CPX_WIDTH-1:0]       cpx_data = fake_iob_out_data;

// Output buffer
// The output buffer need to be asynchronous and cannot ever be overflowed.
// We will ensure this by having a lot of entries
localparam NUM_ASYNC_ENTRIES = 256;

reg [`NOC_DATA_WIDTH-1:0] out_buffer [NUM_ASYNC_ENTRIES-1:0];
reg [NUM_ASYNC_ENTRIES-1:0] out_buffer_val;

reg iob_buffer_val;
reg [2*`NOC_DATA_WIDTH-1:0] iob_buffer_data;

///////////////////////////////////////////////////////////
// write port of the async fifo; runs at chip frequency
///////////////////////////////////////////////////////////
reg [7:0] out_write_index;
reg [7:0] out_write_index_next;

integer i;

always @ (posedge `CHIP.clk_muxed)
begin
    if (!rst_n)
        out_write_index <= 0;
    else
    begin
        out_write_index <= out_write_index_next;
    end

    // write port
    if (!rst_n)
        for (i = 0; i < NUM_ASYNC_ENTRIES; i = i + 1)
        begin
            out_buffer[i] = 0;
            out_buffer_val[i] = 1'b0;
        end
    else
    begin
        if (iob_buffer_val)
        begin
            // no ready; always accepting packet
            out_buffer[out_write_index + 1] = iob_buffer_data[63:0];
            out_buffer[out_write_index] = iob_buffer_data[127:64];
            out_buffer_val[out_write_index] = 1'b1;
            out_buffer_val[out_write_index + 1] = 1'b1;
        end
    end

end

always @ *
begin
    out_write_index_next = iob_buffer_val ? out_write_index + 2 : out_write_index;
end


///////////////////////////////////////////////////////////
// read port of the async fifo; runs at off-chip frequency
///////////////////////////////////////////////////////////
reg [7:0] out_read_index;
reg [7:0] out_read_index_next;

always @ (posedge clk)
begin
    if (!rst_n)
        out_read_index <= 0;
    else
    begin
        out_read_index <= out_read_index_next;
    end

    if (noc_out_rdy && noc_out_val)
    begin
        out_buffer_val[out_read_index] = 1'b0;
    end
end

always @ *
begin
    noc_out_val = out_buffer_val[out_read_index];
    noc_out_data = 0; // Tri: fixes x when out_buffer_counter == 0
    noc_out_data = out_buffer[out_read_index];

    out_read_index_next = (noc_out_rdy && noc_out_val) ? out_read_index + 1 : out_read_index;
end

///////////////////////////////////////////////////////////
// Make out going packets from IOB out data
///////////////////////////////////////////////////////////
reg [63:0] iob_buffer_flit1;
reg [63:0] iob_buffer_flit2;
reg  [`NOC_X_WIDTH-1:0] dest_x;
reg  [`NOC_Y_WIDTH-1:0] dest_y;
always @ *
begin
   iob_buffer_val = fake_iob_out_data[144];
   iob_buffer_flit1 = {14'b0,5'b0, 3'b0, 8'b0,`NOC_FBITS_L1,8'd1, `MSG_TYPE_INTERRUPT,14'b0};
   iob_buffer_flit2 = {fake_iob_out_data[63:16],7'b0,fake_iob_out_data[8:0]};

   // assuming a 8x8 topo
   iob_buffer_flit1[`MSG_DST_X] = dest_x;
   iob_buffer_flit1[`MSG_DST_Y] = dest_y;

   //if (iob_buffer_val)
   //begin
   //   $display("IOB sending to tile X:%d Y:%d", iob_buffer_flit1[`MSG_DST_X], iob_buffer_flit1[`MSG_DST_Y]);
   //   $display("   raw tileid %x", fake_iob_out_data[49:18]);
   // end

   iob_buffer_data = {iob_buffer_flit1, iob_buffer_flit2};
end

always @*
begin
    case (fake_iob_out_data[49:18])
    
32'd0:
begin
    dest_x = `NOC_X_WIDTH'd0;
    dest_y = `NOC_Y_WIDTH'd0;
end

32'd1:
begin
    dest_x = `NOC_X_WIDTH'd1;
    dest_y = `NOC_Y_WIDTH'd0;
end

32'd2:
begin
    dest_x = `NOC_X_WIDTH'd2;
    dest_y = `NOC_Y_WIDTH'd0;
end

32'd3:
begin
    dest_x = `NOC_X_WIDTH'd3;
    dest_y = `NOC_Y_WIDTH'd0;
end

32'd4:
begin
    dest_x = `NOC_X_WIDTH'd4;
    dest_y = `NOC_Y_WIDTH'd0;
end

32'd5:
begin
    dest_x = `NOC_X_WIDTH'd5;
    dest_y = `NOC_Y_WIDTH'd0;
end

32'd6:
begin
    dest_x = `NOC_X_WIDTH'd6;
    dest_y = `NOC_Y_WIDTH'd0;
end

32'd7:
begin
    dest_x = `NOC_X_WIDTH'd7;
    dest_y = `NOC_Y_WIDTH'd0;
end

32'd8:
begin
    dest_x = `NOC_X_WIDTH'd8;
    dest_y = `NOC_Y_WIDTH'd0;
end

32'd9:
begin
    dest_x = `NOC_X_WIDTH'd9;
    dest_y = `NOC_Y_WIDTH'd0;
end

32'd10:
begin
    dest_x = `NOC_X_WIDTH'd10;
    dest_y = `NOC_Y_WIDTH'd0;
end

32'd11:
begin
    dest_x = `NOC_X_WIDTH'd11;
    dest_y = `NOC_Y_WIDTH'd0;
end

32'd12:
begin
    dest_x = `NOC_X_WIDTH'd12;
    dest_y = `NOC_Y_WIDTH'd0;
end

32'd13:
begin
    dest_x = `NOC_X_WIDTH'd13;
    dest_y = `NOC_Y_WIDTH'd0;
end

32'd14:
begin
    dest_x = `NOC_X_WIDTH'd14;
    dest_y = `NOC_Y_WIDTH'd0;
end

32'd15:
begin
    dest_x = `NOC_X_WIDTH'd15;
    dest_y = `NOC_Y_WIDTH'd0;
end

32'd16:
begin
    dest_x = `NOC_X_WIDTH'd16;
    dest_y = `NOC_Y_WIDTH'd0;
end

32'd17:
begin
    dest_x = `NOC_X_WIDTH'd17;
    dest_y = `NOC_Y_WIDTH'd0;
end

32'd18:
begin
    dest_x = `NOC_X_WIDTH'd18;
    dest_y = `NOC_Y_WIDTH'd0;
end

32'd19:
begin
    dest_x = `NOC_X_WIDTH'd19;
    dest_y = `NOC_Y_WIDTH'd0;
end

32'd20:
begin
    dest_x = `NOC_X_WIDTH'd20;
    dest_y = `NOC_Y_WIDTH'd0;
end

32'd21:
begin
    dest_x = `NOC_X_WIDTH'd21;
    dest_y = `NOC_Y_WIDTH'd0;
end

32'd22:
begin
    dest_x = `NOC_X_WIDTH'd22;
    dest_y = `NOC_Y_WIDTH'd0;
end

32'd23:
begin
    dest_x = `NOC_X_WIDTH'd23;
    dest_y = `NOC_Y_WIDTH'd0;
end

32'd24:
begin
    dest_x = `NOC_X_WIDTH'd24;
    dest_y = `NOC_Y_WIDTH'd0;
end

32'd25:
begin
    dest_x = `NOC_X_WIDTH'd25;
    dest_y = `NOC_Y_WIDTH'd0;
end

32'd26:
begin
    dest_x = `NOC_X_WIDTH'd26;
    dest_y = `NOC_Y_WIDTH'd0;
end

32'd27:
begin
    dest_x = `NOC_X_WIDTH'd27;
    dest_y = `NOC_Y_WIDTH'd0;
end

32'd28:
begin
    dest_x = `NOC_X_WIDTH'd28;
    dest_y = `NOC_Y_WIDTH'd0;
end

32'd29:
begin
    dest_x = `NOC_X_WIDTH'd29;
    dest_y = `NOC_Y_WIDTH'd0;
end

32'd30:
begin
    dest_x = `NOC_X_WIDTH'd30;
    dest_y = `NOC_Y_WIDTH'd0;
end

32'd31:
begin
    dest_x = `NOC_X_WIDTH'd31;
    dest_y = `NOC_Y_WIDTH'd0;
end

32'd32:
begin
    dest_x = `NOC_X_WIDTH'd0;
    dest_y = `NOC_Y_WIDTH'd1;
end

32'd33:
begin
    dest_x = `NOC_X_WIDTH'd1;
    dest_y = `NOC_Y_WIDTH'd1;
end

32'd34:
begin
    dest_x = `NOC_X_WIDTH'd2;
    dest_y = `NOC_Y_WIDTH'd1;
end

32'd35:
begin
    dest_x = `NOC_X_WIDTH'd3;
    dest_y = `NOC_Y_WIDTH'd1;
end

32'd36:
begin
    dest_x = `NOC_X_WIDTH'd4;
    dest_y = `NOC_Y_WIDTH'd1;
end

32'd37:
begin
    dest_x = `NOC_X_WIDTH'd5;
    dest_y = `NOC_Y_WIDTH'd1;
end

32'd38:
begin
    dest_x = `NOC_X_WIDTH'd6;
    dest_y = `NOC_Y_WIDTH'd1;
end

32'd39:
begin
    dest_x = `NOC_X_WIDTH'd7;
    dest_y = `NOC_Y_WIDTH'd1;
end

32'd40:
begin
    dest_x = `NOC_X_WIDTH'd8;
    dest_y = `NOC_Y_WIDTH'd1;
end

32'd41:
begin
    dest_x = `NOC_X_WIDTH'd9;
    dest_y = `NOC_Y_WIDTH'd1;
end

32'd42:
begin
    dest_x = `NOC_X_WIDTH'd10;
    dest_y = `NOC_Y_WIDTH'd1;
end

32'd43:
begin
    dest_x = `NOC_X_WIDTH'd11;
    dest_y = `NOC_Y_WIDTH'd1;
end

32'd44:
begin
    dest_x = `NOC_X_WIDTH'd12;
    dest_y = `NOC_Y_WIDTH'd1;
end

32'd45:
begin
    dest_x = `NOC_X_WIDTH'd13;
    dest_y = `NOC_Y_WIDTH'd1;
end

32'd46:
begin
    dest_x = `NOC_X_WIDTH'd14;
    dest_y = `NOC_Y_WIDTH'd1;
end

32'd47:
begin
    dest_x = `NOC_X_WIDTH'd15;
    dest_y = `NOC_Y_WIDTH'd1;
end

32'd48:
begin
    dest_x = `NOC_X_WIDTH'd16;
    dest_y = `NOC_Y_WIDTH'd1;
end

32'd49:
begin
    dest_x = `NOC_X_WIDTH'd17;
    dest_y = `NOC_Y_WIDTH'd1;
end

32'd50:
begin
    dest_x = `NOC_X_WIDTH'd18;
    dest_y = `NOC_Y_WIDTH'd1;
end

32'd51:
begin
    dest_x = `NOC_X_WIDTH'd19;
    dest_y = `NOC_Y_WIDTH'd1;
end

32'd52:
begin
    dest_x = `NOC_X_WIDTH'd20;
    dest_y = `NOC_Y_WIDTH'd1;
end

32'd53:
begin
    dest_x = `NOC_X_WIDTH'd21;
    dest_y = `NOC_Y_WIDTH'd1;
end

32'd54:
begin
    dest_x = `NOC_X_WIDTH'd22;
    dest_y = `NOC_Y_WIDTH'd1;
end

32'd55:
begin
    dest_x = `NOC_X_WIDTH'd23;
    dest_y = `NOC_Y_WIDTH'd1;
end

32'd56:
begin
    dest_x = `NOC_X_WIDTH'd24;
    dest_y = `NOC_Y_WIDTH'd1;
end

32'd57:
begin
    dest_x = `NOC_X_WIDTH'd25;
    dest_y = `NOC_Y_WIDTH'd1;
end

32'd58:
begin
    dest_x = `NOC_X_WIDTH'd26;
    dest_y = `NOC_Y_WIDTH'd1;
end

32'd59:
begin
    dest_x = `NOC_X_WIDTH'd27;
    dest_y = `NOC_Y_WIDTH'd1;
end

32'd60:
begin
    dest_x = `NOC_X_WIDTH'd28;
    dest_y = `NOC_Y_WIDTH'd1;
end

32'd61:
begin
    dest_x = `NOC_X_WIDTH'd29;
    dest_y = `NOC_Y_WIDTH'd1;
end

32'd62:
begin
    dest_x = `NOC_X_WIDTH'd30;
    dest_y = `NOC_Y_WIDTH'd1;
end

32'd63:
begin
    dest_x = `NOC_X_WIDTH'd31;
    dest_y = `NOC_Y_WIDTH'd1;
end

32'd64:
begin
    dest_x = `NOC_X_WIDTH'd0;
    dest_y = `NOC_Y_WIDTH'd2;
end

32'd65:
begin
    dest_x = `NOC_X_WIDTH'd1;
    dest_y = `NOC_Y_WIDTH'd2;
end

32'd66:
begin
    dest_x = `NOC_X_WIDTH'd2;
    dest_y = `NOC_Y_WIDTH'd2;
end

32'd67:
begin
    dest_x = `NOC_X_WIDTH'd3;
    dest_y = `NOC_Y_WIDTH'd2;
end

32'd68:
begin
    dest_x = `NOC_X_WIDTH'd4;
    dest_y = `NOC_Y_WIDTH'd2;
end

32'd69:
begin
    dest_x = `NOC_X_WIDTH'd5;
    dest_y = `NOC_Y_WIDTH'd2;
end

32'd70:
begin
    dest_x = `NOC_X_WIDTH'd6;
    dest_y = `NOC_Y_WIDTH'd2;
end

32'd71:
begin
    dest_x = `NOC_X_WIDTH'd7;
    dest_y = `NOC_Y_WIDTH'd2;
end

32'd72:
begin
    dest_x = `NOC_X_WIDTH'd8;
    dest_y = `NOC_Y_WIDTH'd2;
end

32'd73:
begin
    dest_x = `NOC_X_WIDTH'd9;
    dest_y = `NOC_Y_WIDTH'd2;
end

32'd74:
begin
    dest_x = `NOC_X_WIDTH'd10;
    dest_y = `NOC_Y_WIDTH'd2;
end

32'd75:
begin
    dest_x = `NOC_X_WIDTH'd11;
    dest_y = `NOC_Y_WIDTH'd2;
end

32'd76:
begin
    dest_x = `NOC_X_WIDTH'd12;
    dest_y = `NOC_Y_WIDTH'd2;
end

32'd77:
begin
    dest_x = `NOC_X_WIDTH'd13;
    dest_y = `NOC_Y_WIDTH'd2;
end

32'd78:
begin
    dest_x = `NOC_X_WIDTH'd14;
    dest_y = `NOC_Y_WIDTH'd2;
end

32'd79:
begin
    dest_x = `NOC_X_WIDTH'd15;
    dest_y = `NOC_Y_WIDTH'd2;
end

32'd80:
begin
    dest_x = `NOC_X_WIDTH'd16;
    dest_y = `NOC_Y_WIDTH'd2;
end

32'd81:
begin
    dest_x = `NOC_X_WIDTH'd17;
    dest_y = `NOC_Y_WIDTH'd2;
end

32'd82:
begin
    dest_x = `NOC_X_WIDTH'd18;
    dest_y = `NOC_Y_WIDTH'd2;
end

32'd83:
begin
    dest_x = `NOC_X_WIDTH'd19;
    dest_y = `NOC_Y_WIDTH'd2;
end

32'd84:
begin
    dest_x = `NOC_X_WIDTH'd20;
    dest_y = `NOC_Y_WIDTH'd2;
end

32'd85:
begin
    dest_x = `NOC_X_WIDTH'd21;
    dest_y = `NOC_Y_WIDTH'd2;
end

32'd86:
begin
    dest_x = `NOC_X_WIDTH'd22;
    dest_y = `NOC_Y_WIDTH'd2;
end

32'd87:
begin
    dest_x = `NOC_X_WIDTH'd23;
    dest_y = `NOC_Y_WIDTH'd2;
end

32'd88:
begin
    dest_x = `NOC_X_WIDTH'd24;
    dest_y = `NOC_Y_WIDTH'd2;
end

32'd89:
begin
    dest_x = `NOC_X_WIDTH'd25;
    dest_y = `NOC_Y_WIDTH'd2;
end

32'd90:
begin
    dest_x = `NOC_X_WIDTH'd26;
    dest_y = `NOC_Y_WIDTH'd2;
end

32'd91:
begin
    dest_x = `NOC_X_WIDTH'd27;
    dest_y = `NOC_Y_WIDTH'd2;
end

32'd92:
begin
    dest_x = `NOC_X_WIDTH'd28;
    dest_y = `NOC_Y_WIDTH'd2;
end

32'd93:
begin
    dest_x = `NOC_X_WIDTH'd29;
    dest_y = `NOC_Y_WIDTH'd2;
end

32'd94:
begin
    dest_x = `NOC_X_WIDTH'd30;
    dest_y = `NOC_Y_WIDTH'd2;
end

32'd95:
begin
    dest_x = `NOC_X_WIDTH'd31;
    dest_y = `NOC_Y_WIDTH'd2;
end

32'd96:
begin
    dest_x = `NOC_X_WIDTH'd0;
    dest_y = `NOC_Y_WIDTH'd3;
end

32'd97:
begin
    dest_x = `NOC_X_WIDTH'd1;
    dest_y = `NOC_Y_WIDTH'd3;
end

32'd98:
begin
    dest_x = `NOC_X_WIDTH'd2;
    dest_y = `NOC_Y_WIDTH'd3;
end

32'd99:
begin
    dest_x = `NOC_X_WIDTH'd3;
    dest_y = `NOC_Y_WIDTH'd3;
end

32'd100:
begin
    dest_x = `NOC_X_WIDTH'd4;
    dest_y = `NOC_Y_WIDTH'd3;
end

32'd101:
begin
    dest_x = `NOC_X_WIDTH'd5;
    dest_y = `NOC_Y_WIDTH'd3;
end

32'd102:
begin
    dest_x = `NOC_X_WIDTH'd6;
    dest_y = `NOC_Y_WIDTH'd3;
end

32'd103:
begin
    dest_x = `NOC_X_WIDTH'd7;
    dest_y = `NOC_Y_WIDTH'd3;
end

32'd104:
begin
    dest_x = `NOC_X_WIDTH'd8;
    dest_y = `NOC_Y_WIDTH'd3;
end

32'd105:
begin
    dest_x = `NOC_X_WIDTH'd9;
    dest_y = `NOC_Y_WIDTH'd3;
end

32'd106:
begin
    dest_x = `NOC_X_WIDTH'd10;
    dest_y = `NOC_Y_WIDTH'd3;
end

32'd107:
begin
    dest_x = `NOC_X_WIDTH'd11;
    dest_y = `NOC_Y_WIDTH'd3;
end

32'd108:
begin
    dest_x = `NOC_X_WIDTH'd12;
    dest_y = `NOC_Y_WIDTH'd3;
end

32'd109:
begin
    dest_x = `NOC_X_WIDTH'd13;
    dest_y = `NOC_Y_WIDTH'd3;
end

32'd110:
begin
    dest_x = `NOC_X_WIDTH'd14;
    dest_y = `NOC_Y_WIDTH'd3;
end

32'd111:
begin
    dest_x = `NOC_X_WIDTH'd15;
    dest_y = `NOC_Y_WIDTH'd3;
end

32'd112:
begin
    dest_x = `NOC_X_WIDTH'd16;
    dest_y = `NOC_Y_WIDTH'd3;
end

32'd113:
begin
    dest_x = `NOC_X_WIDTH'd17;
    dest_y = `NOC_Y_WIDTH'd3;
end

32'd114:
begin
    dest_x = `NOC_X_WIDTH'd18;
    dest_y = `NOC_Y_WIDTH'd3;
end

32'd115:
begin
    dest_x = `NOC_X_WIDTH'd19;
    dest_y = `NOC_Y_WIDTH'd3;
end

32'd116:
begin
    dest_x = `NOC_X_WIDTH'd20;
    dest_y = `NOC_Y_WIDTH'd3;
end

32'd117:
begin
    dest_x = `NOC_X_WIDTH'd21;
    dest_y = `NOC_Y_WIDTH'd3;
end

32'd118:
begin
    dest_x = `NOC_X_WIDTH'd22;
    dest_y = `NOC_Y_WIDTH'd3;
end

32'd119:
begin
    dest_x = `NOC_X_WIDTH'd23;
    dest_y = `NOC_Y_WIDTH'd3;
end

32'd120:
begin
    dest_x = `NOC_X_WIDTH'd24;
    dest_y = `NOC_Y_WIDTH'd3;
end

32'd121:
begin
    dest_x = `NOC_X_WIDTH'd25;
    dest_y = `NOC_Y_WIDTH'd3;
end

32'd122:
begin
    dest_x = `NOC_X_WIDTH'd26;
    dest_y = `NOC_Y_WIDTH'd3;
end

32'd123:
begin
    dest_x = `NOC_X_WIDTH'd27;
    dest_y = `NOC_Y_WIDTH'd3;
end

32'd124:
begin
    dest_x = `NOC_X_WIDTH'd28;
    dest_y = `NOC_Y_WIDTH'd3;
end

32'd125:
begin
    dest_x = `NOC_X_WIDTH'd29;
    dest_y = `NOC_Y_WIDTH'd3;
end

32'd126:
begin
    dest_x = `NOC_X_WIDTH'd30;
    dest_y = `NOC_Y_WIDTH'd3;
end

32'd127:
begin
    dest_x = `NOC_X_WIDTH'd31;
    dest_y = `NOC_Y_WIDTH'd3;
end

32'd128:
begin
    dest_x = `NOC_X_WIDTH'd0;
    dest_y = `NOC_Y_WIDTH'd4;
end

32'd129:
begin
    dest_x = `NOC_X_WIDTH'd1;
    dest_y = `NOC_Y_WIDTH'd4;
end

32'd130:
begin
    dest_x = `NOC_X_WIDTH'd2;
    dest_y = `NOC_Y_WIDTH'd4;
end

32'd131:
begin
    dest_x = `NOC_X_WIDTH'd3;
    dest_y = `NOC_Y_WIDTH'd4;
end

32'd132:
begin
    dest_x = `NOC_X_WIDTH'd4;
    dest_y = `NOC_Y_WIDTH'd4;
end

32'd133:
begin
    dest_x = `NOC_X_WIDTH'd5;
    dest_y = `NOC_Y_WIDTH'd4;
end

32'd134:
begin
    dest_x = `NOC_X_WIDTH'd6;
    dest_y = `NOC_Y_WIDTH'd4;
end

32'd135:
begin
    dest_x = `NOC_X_WIDTH'd7;
    dest_y = `NOC_Y_WIDTH'd4;
end

32'd136:
begin
    dest_x = `NOC_X_WIDTH'd8;
    dest_y = `NOC_Y_WIDTH'd4;
end

32'd137:
begin
    dest_x = `NOC_X_WIDTH'd9;
    dest_y = `NOC_Y_WIDTH'd4;
end

32'd138:
begin
    dest_x = `NOC_X_WIDTH'd10;
    dest_y = `NOC_Y_WIDTH'd4;
end

32'd139:
begin
    dest_x = `NOC_X_WIDTH'd11;
    dest_y = `NOC_Y_WIDTH'd4;
end

32'd140:
begin
    dest_x = `NOC_X_WIDTH'd12;
    dest_y = `NOC_Y_WIDTH'd4;
end

32'd141:
begin
    dest_x = `NOC_X_WIDTH'd13;
    dest_y = `NOC_Y_WIDTH'd4;
end

32'd142:
begin
    dest_x = `NOC_X_WIDTH'd14;
    dest_y = `NOC_Y_WIDTH'd4;
end

32'd143:
begin
    dest_x = `NOC_X_WIDTH'd15;
    dest_y = `NOC_Y_WIDTH'd4;
end

32'd144:
begin
    dest_x = `NOC_X_WIDTH'd16;
    dest_y = `NOC_Y_WIDTH'd4;
end

32'd145:
begin
    dest_x = `NOC_X_WIDTH'd17;
    dest_y = `NOC_Y_WIDTH'd4;
end

32'd146:
begin
    dest_x = `NOC_X_WIDTH'd18;
    dest_y = `NOC_Y_WIDTH'd4;
end

32'd147:
begin
    dest_x = `NOC_X_WIDTH'd19;
    dest_y = `NOC_Y_WIDTH'd4;
end

32'd148:
begin
    dest_x = `NOC_X_WIDTH'd20;
    dest_y = `NOC_Y_WIDTH'd4;
end

32'd149:
begin
    dest_x = `NOC_X_WIDTH'd21;
    dest_y = `NOC_Y_WIDTH'd4;
end

32'd150:
begin
    dest_x = `NOC_X_WIDTH'd22;
    dest_y = `NOC_Y_WIDTH'd4;
end

32'd151:
begin
    dest_x = `NOC_X_WIDTH'd23;
    dest_y = `NOC_Y_WIDTH'd4;
end

32'd152:
begin
    dest_x = `NOC_X_WIDTH'd24;
    dest_y = `NOC_Y_WIDTH'd4;
end

32'd153:
begin
    dest_x = `NOC_X_WIDTH'd25;
    dest_y = `NOC_Y_WIDTH'd4;
end

32'd154:
begin
    dest_x = `NOC_X_WIDTH'd26;
    dest_y = `NOC_Y_WIDTH'd4;
end

32'd155:
begin
    dest_x = `NOC_X_WIDTH'd27;
    dest_y = `NOC_Y_WIDTH'd4;
end

32'd156:
begin
    dest_x = `NOC_X_WIDTH'd28;
    dest_y = `NOC_Y_WIDTH'd4;
end

32'd157:
begin
    dest_x = `NOC_X_WIDTH'd29;
    dest_y = `NOC_Y_WIDTH'd4;
end

32'd158:
begin
    dest_x = `NOC_X_WIDTH'd30;
    dest_y = `NOC_Y_WIDTH'd4;
end

32'd159:
begin
    dest_x = `NOC_X_WIDTH'd31;
    dest_y = `NOC_Y_WIDTH'd4;
end

32'd160:
begin
    dest_x = `NOC_X_WIDTH'd0;
    dest_y = `NOC_Y_WIDTH'd5;
end

32'd161:
begin
    dest_x = `NOC_X_WIDTH'd1;
    dest_y = `NOC_Y_WIDTH'd5;
end

32'd162:
begin
    dest_x = `NOC_X_WIDTH'd2;
    dest_y = `NOC_Y_WIDTH'd5;
end

32'd163:
begin
    dest_x = `NOC_X_WIDTH'd3;
    dest_y = `NOC_Y_WIDTH'd5;
end

32'd164:
begin
    dest_x = `NOC_X_WIDTH'd4;
    dest_y = `NOC_Y_WIDTH'd5;
end

32'd165:
begin
    dest_x = `NOC_X_WIDTH'd5;
    dest_y = `NOC_Y_WIDTH'd5;
end

32'd166:
begin
    dest_x = `NOC_X_WIDTH'd6;
    dest_y = `NOC_Y_WIDTH'd5;
end

32'd167:
begin
    dest_x = `NOC_X_WIDTH'd7;
    dest_y = `NOC_Y_WIDTH'd5;
end

32'd168:
begin
    dest_x = `NOC_X_WIDTH'd8;
    dest_y = `NOC_Y_WIDTH'd5;
end

32'd169:
begin
    dest_x = `NOC_X_WIDTH'd9;
    dest_y = `NOC_Y_WIDTH'd5;
end

32'd170:
begin
    dest_x = `NOC_X_WIDTH'd10;
    dest_y = `NOC_Y_WIDTH'd5;
end

32'd171:
begin
    dest_x = `NOC_X_WIDTH'd11;
    dest_y = `NOC_Y_WIDTH'd5;
end

32'd172:
begin
    dest_x = `NOC_X_WIDTH'd12;
    dest_y = `NOC_Y_WIDTH'd5;
end

32'd173:
begin
    dest_x = `NOC_X_WIDTH'd13;
    dest_y = `NOC_Y_WIDTH'd5;
end

32'd174:
begin
    dest_x = `NOC_X_WIDTH'd14;
    dest_y = `NOC_Y_WIDTH'd5;
end

32'd175:
begin
    dest_x = `NOC_X_WIDTH'd15;
    dest_y = `NOC_Y_WIDTH'd5;
end

32'd176:
begin
    dest_x = `NOC_X_WIDTH'd16;
    dest_y = `NOC_Y_WIDTH'd5;
end

32'd177:
begin
    dest_x = `NOC_X_WIDTH'd17;
    dest_y = `NOC_Y_WIDTH'd5;
end

32'd178:
begin
    dest_x = `NOC_X_WIDTH'd18;
    dest_y = `NOC_Y_WIDTH'd5;
end

32'd179:
begin
    dest_x = `NOC_X_WIDTH'd19;
    dest_y = `NOC_Y_WIDTH'd5;
end

32'd180:
begin
    dest_x = `NOC_X_WIDTH'd20;
    dest_y = `NOC_Y_WIDTH'd5;
end

32'd181:
begin
    dest_x = `NOC_X_WIDTH'd21;
    dest_y = `NOC_Y_WIDTH'd5;
end

32'd182:
begin
    dest_x = `NOC_X_WIDTH'd22;
    dest_y = `NOC_Y_WIDTH'd5;
end

32'd183:
begin
    dest_x = `NOC_X_WIDTH'd23;
    dest_y = `NOC_Y_WIDTH'd5;
end

32'd184:
begin
    dest_x = `NOC_X_WIDTH'd24;
    dest_y = `NOC_Y_WIDTH'd5;
end

32'd185:
begin
    dest_x = `NOC_X_WIDTH'd25;
    dest_y = `NOC_Y_WIDTH'd5;
end

32'd186:
begin
    dest_x = `NOC_X_WIDTH'd26;
    dest_y = `NOC_Y_WIDTH'd5;
end

32'd187:
begin
    dest_x = `NOC_X_WIDTH'd27;
    dest_y = `NOC_Y_WIDTH'd5;
end

32'd188:
begin
    dest_x = `NOC_X_WIDTH'd28;
    dest_y = `NOC_Y_WIDTH'd5;
end

32'd189:
begin
    dest_x = `NOC_X_WIDTH'd29;
    dest_y = `NOC_Y_WIDTH'd5;
end

32'd190:
begin
    dest_x = `NOC_X_WIDTH'd30;
    dest_y = `NOC_Y_WIDTH'd5;
end

32'd191:
begin
    dest_x = `NOC_X_WIDTH'd31;
    dest_y = `NOC_Y_WIDTH'd5;
end

32'd192:
begin
    dest_x = `NOC_X_WIDTH'd0;
    dest_y = `NOC_Y_WIDTH'd6;
end

32'd193:
begin
    dest_x = `NOC_X_WIDTH'd1;
    dest_y = `NOC_Y_WIDTH'd6;
end

32'd194:
begin
    dest_x = `NOC_X_WIDTH'd2;
    dest_y = `NOC_Y_WIDTH'd6;
end

32'd195:
begin
    dest_x = `NOC_X_WIDTH'd3;
    dest_y = `NOC_Y_WIDTH'd6;
end

32'd196:
begin
    dest_x = `NOC_X_WIDTH'd4;
    dest_y = `NOC_Y_WIDTH'd6;
end

32'd197:
begin
    dest_x = `NOC_X_WIDTH'd5;
    dest_y = `NOC_Y_WIDTH'd6;
end

32'd198:
begin
    dest_x = `NOC_X_WIDTH'd6;
    dest_y = `NOC_Y_WIDTH'd6;
end

32'd199:
begin
    dest_x = `NOC_X_WIDTH'd7;
    dest_y = `NOC_Y_WIDTH'd6;
end

32'd200:
begin
    dest_x = `NOC_X_WIDTH'd8;
    dest_y = `NOC_Y_WIDTH'd6;
end

32'd201:
begin
    dest_x = `NOC_X_WIDTH'd9;
    dest_y = `NOC_Y_WIDTH'd6;
end

32'd202:
begin
    dest_x = `NOC_X_WIDTH'd10;
    dest_y = `NOC_Y_WIDTH'd6;
end

32'd203:
begin
    dest_x = `NOC_X_WIDTH'd11;
    dest_y = `NOC_Y_WIDTH'd6;
end

32'd204:
begin
    dest_x = `NOC_X_WIDTH'd12;
    dest_y = `NOC_Y_WIDTH'd6;
end

32'd205:
begin
    dest_x = `NOC_X_WIDTH'd13;
    dest_y = `NOC_Y_WIDTH'd6;
end

32'd206:
begin
    dest_x = `NOC_X_WIDTH'd14;
    dest_y = `NOC_Y_WIDTH'd6;
end

32'd207:
begin
    dest_x = `NOC_X_WIDTH'd15;
    dest_y = `NOC_Y_WIDTH'd6;
end

32'd208:
begin
    dest_x = `NOC_X_WIDTH'd16;
    dest_y = `NOC_Y_WIDTH'd6;
end

32'd209:
begin
    dest_x = `NOC_X_WIDTH'd17;
    dest_y = `NOC_Y_WIDTH'd6;
end

32'd210:
begin
    dest_x = `NOC_X_WIDTH'd18;
    dest_y = `NOC_Y_WIDTH'd6;
end

32'd211:
begin
    dest_x = `NOC_X_WIDTH'd19;
    dest_y = `NOC_Y_WIDTH'd6;
end

32'd212:
begin
    dest_x = `NOC_X_WIDTH'd20;
    dest_y = `NOC_Y_WIDTH'd6;
end

32'd213:
begin
    dest_x = `NOC_X_WIDTH'd21;
    dest_y = `NOC_Y_WIDTH'd6;
end

32'd214:
begin
    dest_x = `NOC_X_WIDTH'd22;
    dest_y = `NOC_Y_WIDTH'd6;
end

32'd215:
begin
    dest_x = `NOC_X_WIDTH'd23;
    dest_y = `NOC_Y_WIDTH'd6;
end

32'd216:
begin
    dest_x = `NOC_X_WIDTH'd24;
    dest_y = `NOC_Y_WIDTH'd6;
end

32'd217:
begin
    dest_x = `NOC_X_WIDTH'd25;
    dest_y = `NOC_Y_WIDTH'd6;
end

32'd218:
begin
    dest_x = `NOC_X_WIDTH'd26;
    dest_y = `NOC_Y_WIDTH'd6;
end

32'd219:
begin
    dest_x = `NOC_X_WIDTH'd27;
    dest_y = `NOC_Y_WIDTH'd6;
end

32'd220:
begin
    dest_x = `NOC_X_WIDTH'd28;
    dest_y = `NOC_Y_WIDTH'd6;
end

32'd221:
begin
    dest_x = `NOC_X_WIDTH'd29;
    dest_y = `NOC_Y_WIDTH'd6;
end

32'd222:
begin
    dest_x = `NOC_X_WIDTH'd30;
    dest_y = `NOC_Y_WIDTH'd6;
end

32'd223:
begin
    dest_x = `NOC_X_WIDTH'd31;
    dest_y = `NOC_Y_WIDTH'd6;
end

32'd224:
begin
    dest_x = `NOC_X_WIDTH'd0;
    dest_y = `NOC_Y_WIDTH'd7;
end

32'd225:
begin
    dest_x = `NOC_X_WIDTH'd1;
    dest_y = `NOC_Y_WIDTH'd7;
end

32'd226:
begin
    dest_x = `NOC_X_WIDTH'd2;
    dest_y = `NOC_Y_WIDTH'd7;
end

32'd227:
begin
    dest_x = `NOC_X_WIDTH'd3;
    dest_y = `NOC_Y_WIDTH'd7;
end

32'd228:
begin
    dest_x = `NOC_X_WIDTH'd4;
    dest_y = `NOC_Y_WIDTH'd7;
end

32'd229:
begin
    dest_x = `NOC_X_WIDTH'd5;
    dest_y = `NOC_Y_WIDTH'd7;
end

32'd230:
begin
    dest_x = `NOC_X_WIDTH'd6;
    dest_y = `NOC_Y_WIDTH'd7;
end

32'd231:
begin
    dest_x = `NOC_X_WIDTH'd7;
    dest_y = `NOC_Y_WIDTH'd7;
end

32'd232:
begin
    dest_x = `NOC_X_WIDTH'd8;
    dest_y = `NOC_Y_WIDTH'd7;
end

32'd233:
begin
    dest_x = `NOC_X_WIDTH'd9;
    dest_y = `NOC_Y_WIDTH'd7;
end

32'd234:
begin
    dest_x = `NOC_X_WIDTH'd10;
    dest_y = `NOC_Y_WIDTH'd7;
end

32'd235:
begin
    dest_x = `NOC_X_WIDTH'd11;
    dest_y = `NOC_Y_WIDTH'd7;
end

32'd236:
begin
    dest_x = `NOC_X_WIDTH'd12;
    dest_y = `NOC_Y_WIDTH'd7;
end

32'd237:
begin
    dest_x = `NOC_X_WIDTH'd13;
    dest_y = `NOC_Y_WIDTH'd7;
end

32'd238:
begin
    dest_x = `NOC_X_WIDTH'd14;
    dest_y = `NOC_Y_WIDTH'd7;
end

32'd239:
begin
    dest_x = `NOC_X_WIDTH'd15;
    dest_y = `NOC_Y_WIDTH'd7;
end

32'd240:
begin
    dest_x = `NOC_X_WIDTH'd16;
    dest_y = `NOC_Y_WIDTH'd7;
end

32'd241:
begin
    dest_x = `NOC_X_WIDTH'd17;
    dest_y = `NOC_Y_WIDTH'd7;
end

32'd242:
begin
    dest_x = `NOC_X_WIDTH'd18;
    dest_y = `NOC_Y_WIDTH'd7;
end

32'd243:
begin
    dest_x = `NOC_X_WIDTH'd19;
    dest_y = `NOC_Y_WIDTH'd7;
end

32'd244:
begin
    dest_x = `NOC_X_WIDTH'd20;
    dest_y = `NOC_Y_WIDTH'd7;
end

32'd245:
begin
    dest_x = `NOC_X_WIDTH'd21;
    dest_y = `NOC_Y_WIDTH'd7;
end

32'd246:
begin
    dest_x = `NOC_X_WIDTH'd22;
    dest_y = `NOC_Y_WIDTH'd7;
end

32'd247:
begin
    dest_x = `NOC_X_WIDTH'd23;
    dest_y = `NOC_Y_WIDTH'd7;
end

32'd248:
begin
    dest_x = `NOC_X_WIDTH'd24;
    dest_y = `NOC_Y_WIDTH'd7;
end

32'd249:
begin
    dest_x = `NOC_X_WIDTH'd25;
    dest_y = `NOC_Y_WIDTH'd7;
end

32'd250:
begin
    dest_x = `NOC_X_WIDTH'd26;
    dest_y = `NOC_Y_WIDTH'd7;
end

32'd251:
begin
    dest_x = `NOC_X_WIDTH'd27;
    dest_y = `NOC_Y_WIDTH'd7;
end

32'd252:
begin
    dest_x = `NOC_X_WIDTH'd28;
    dest_y = `NOC_Y_WIDTH'd7;
end

32'd253:
begin
    dest_x = `NOC_X_WIDTH'd29;
    dest_y = `NOC_Y_WIDTH'd7;
end

32'd254:
begin
    dest_x = `NOC_X_WIDTH'd30;
    dest_y = `NOC_Y_WIDTH'd7;
end

32'd255:
begin
    dest_x = `NOC_X_WIDTH'd31;
    dest_y = `NOC_Y_WIDTH'd7;
end

32'd256:
begin
    dest_x = `NOC_X_WIDTH'd0;
    dest_y = `NOC_Y_WIDTH'd8;
end

32'd257:
begin
    dest_x = `NOC_X_WIDTH'd1;
    dest_y = `NOC_Y_WIDTH'd8;
end

32'd258:
begin
    dest_x = `NOC_X_WIDTH'd2;
    dest_y = `NOC_Y_WIDTH'd8;
end

32'd259:
begin
    dest_x = `NOC_X_WIDTH'd3;
    dest_y = `NOC_Y_WIDTH'd8;
end

32'd260:
begin
    dest_x = `NOC_X_WIDTH'd4;
    dest_y = `NOC_Y_WIDTH'd8;
end

32'd261:
begin
    dest_x = `NOC_X_WIDTH'd5;
    dest_y = `NOC_Y_WIDTH'd8;
end

32'd262:
begin
    dest_x = `NOC_X_WIDTH'd6;
    dest_y = `NOC_Y_WIDTH'd8;
end

32'd263:
begin
    dest_x = `NOC_X_WIDTH'd7;
    dest_y = `NOC_Y_WIDTH'd8;
end

32'd264:
begin
    dest_x = `NOC_X_WIDTH'd8;
    dest_y = `NOC_Y_WIDTH'd8;
end

32'd265:
begin
    dest_x = `NOC_X_WIDTH'd9;
    dest_y = `NOC_Y_WIDTH'd8;
end

32'd266:
begin
    dest_x = `NOC_X_WIDTH'd10;
    dest_y = `NOC_Y_WIDTH'd8;
end

32'd267:
begin
    dest_x = `NOC_X_WIDTH'd11;
    dest_y = `NOC_Y_WIDTH'd8;
end

32'd268:
begin
    dest_x = `NOC_X_WIDTH'd12;
    dest_y = `NOC_Y_WIDTH'd8;
end

32'd269:
begin
    dest_x = `NOC_X_WIDTH'd13;
    dest_y = `NOC_Y_WIDTH'd8;
end

32'd270:
begin
    dest_x = `NOC_X_WIDTH'd14;
    dest_y = `NOC_Y_WIDTH'd8;
end

32'd271:
begin
    dest_x = `NOC_X_WIDTH'd15;
    dest_y = `NOC_Y_WIDTH'd8;
end

32'd272:
begin
    dest_x = `NOC_X_WIDTH'd16;
    dest_y = `NOC_Y_WIDTH'd8;
end

32'd273:
begin
    dest_x = `NOC_X_WIDTH'd17;
    dest_y = `NOC_Y_WIDTH'd8;
end

32'd274:
begin
    dest_x = `NOC_X_WIDTH'd18;
    dest_y = `NOC_Y_WIDTH'd8;
end

32'd275:
begin
    dest_x = `NOC_X_WIDTH'd19;
    dest_y = `NOC_Y_WIDTH'd8;
end

32'd276:
begin
    dest_x = `NOC_X_WIDTH'd20;
    dest_y = `NOC_Y_WIDTH'd8;
end

32'd277:
begin
    dest_x = `NOC_X_WIDTH'd21;
    dest_y = `NOC_Y_WIDTH'd8;
end

32'd278:
begin
    dest_x = `NOC_X_WIDTH'd22;
    dest_y = `NOC_Y_WIDTH'd8;
end

32'd279:
begin
    dest_x = `NOC_X_WIDTH'd23;
    dest_y = `NOC_Y_WIDTH'd8;
end

32'd280:
begin
    dest_x = `NOC_X_WIDTH'd24;
    dest_y = `NOC_Y_WIDTH'd8;
end

32'd281:
begin
    dest_x = `NOC_X_WIDTH'd25;
    dest_y = `NOC_Y_WIDTH'd8;
end

32'd282:
begin
    dest_x = `NOC_X_WIDTH'd26;
    dest_y = `NOC_Y_WIDTH'd8;
end

32'd283:
begin
    dest_x = `NOC_X_WIDTH'd27;
    dest_y = `NOC_Y_WIDTH'd8;
end

32'd284:
begin
    dest_x = `NOC_X_WIDTH'd28;
    dest_y = `NOC_Y_WIDTH'd8;
end

32'd285:
begin
    dest_x = `NOC_X_WIDTH'd29;
    dest_y = `NOC_Y_WIDTH'd8;
end

32'd286:
begin
    dest_x = `NOC_X_WIDTH'd30;
    dest_y = `NOC_Y_WIDTH'd8;
end

32'd287:
begin
    dest_x = `NOC_X_WIDTH'd31;
    dest_y = `NOC_Y_WIDTH'd8;
end

32'd288:
begin
    dest_x = `NOC_X_WIDTH'd0;
    dest_y = `NOC_Y_WIDTH'd9;
end

32'd289:
begin
    dest_x = `NOC_X_WIDTH'd1;
    dest_y = `NOC_Y_WIDTH'd9;
end

32'd290:
begin
    dest_x = `NOC_X_WIDTH'd2;
    dest_y = `NOC_Y_WIDTH'd9;
end

32'd291:
begin
    dest_x = `NOC_X_WIDTH'd3;
    dest_y = `NOC_Y_WIDTH'd9;
end

32'd292:
begin
    dest_x = `NOC_X_WIDTH'd4;
    dest_y = `NOC_Y_WIDTH'd9;
end

32'd293:
begin
    dest_x = `NOC_X_WIDTH'd5;
    dest_y = `NOC_Y_WIDTH'd9;
end

32'd294:
begin
    dest_x = `NOC_X_WIDTH'd6;
    dest_y = `NOC_Y_WIDTH'd9;
end

32'd295:
begin
    dest_x = `NOC_X_WIDTH'd7;
    dest_y = `NOC_Y_WIDTH'd9;
end

32'd296:
begin
    dest_x = `NOC_X_WIDTH'd8;
    dest_y = `NOC_Y_WIDTH'd9;
end

32'd297:
begin
    dest_x = `NOC_X_WIDTH'd9;
    dest_y = `NOC_Y_WIDTH'd9;
end

32'd298:
begin
    dest_x = `NOC_X_WIDTH'd10;
    dest_y = `NOC_Y_WIDTH'd9;
end

32'd299:
begin
    dest_x = `NOC_X_WIDTH'd11;
    dest_y = `NOC_Y_WIDTH'd9;
end

32'd300:
begin
    dest_x = `NOC_X_WIDTH'd12;
    dest_y = `NOC_Y_WIDTH'd9;
end

32'd301:
begin
    dest_x = `NOC_X_WIDTH'd13;
    dest_y = `NOC_Y_WIDTH'd9;
end

32'd302:
begin
    dest_x = `NOC_X_WIDTH'd14;
    dest_y = `NOC_Y_WIDTH'd9;
end

32'd303:
begin
    dest_x = `NOC_X_WIDTH'd15;
    dest_y = `NOC_Y_WIDTH'd9;
end

32'd304:
begin
    dest_x = `NOC_X_WIDTH'd16;
    dest_y = `NOC_Y_WIDTH'd9;
end

32'd305:
begin
    dest_x = `NOC_X_WIDTH'd17;
    dest_y = `NOC_Y_WIDTH'd9;
end

32'd306:
begin
    dest_x = `NOC_X_WIDTH'd18;
    dest_y = `NOC_Y_WIDTH'd9;
end

32'd307:
begin
    dest_x = `NOC_X_WIDTH'd19;
    dest_y = `NOC_Y_WIDTH'd9;
end

32'd308:
begin
    dest_x = `NOC_X_WIDTH'd20;
    dest_y = `NOC_Y_WIDTH'd9;
end

32'd309:
begin
    dest_x = `NOC_X_WIDTH'd21;
    dest_y = `NOC_Y_WIDTH'd9;
end

32'd310:
begin
    dest_x = `NOC_X_WIDTH'd22;
    dest_y = `NOC_Y_WIDTH'd9;
end

32'd311:
begin
    dest_x = `NOC_X_WIDTH'd23;
    dest_y = `NOC_Y_WIDTH'd9;
end

32'd312:
begin
    dest_x = `NOC_X_WIDTH'd24;
    dest_y = `NOC_Y_WIDTH'd9;
end

32'd313:
begin
    dest_x = `NOC_X_WIDTH'd25;
    dest_y = `NOC_Y_WIDTH'd9;
end

32'd314:
begin
    dest_x = `NOC_X_WIDTH'd26;
    dest_y = `NOC_Y_WIDTH'd9;
end

32'd315:
begin
    dest_x = `NOC_X_WIDTH'd27;
    dest_y = `NOC_Y_WIDTH'd9;
end

32'd316:
begin
    dest_x = `NOC_X_WIDTH'd28;
    dest_y = `NOC_Y_WIDTH'd9;
end

32'd317:
begin
    dest_x = `NOC_X_WIDTH'd29;
    dest_y = `NOC_Y_WIDTH'd9;
end

32'd318:
begin
    dest_x = `NOC_X_WIDTH'd30;
    dest_y = `NOC_Y_WIDTH'd9;
end

32'd319:
begin
    dest_x = `NOC_X_WIDTH'd31;
    dest_y = `NOC_Y_WIDTH'd9;
end

32'd320:
begin
    dest_x = `NOC_X_WIDTH'd0;
    dest_y = `NOC_Y_WIDTH'd10;
end

32'd321:
begin
    dest_x = `NOC_X_WIDTH'd1;
    dest_y = `NOC_Y_WIDTH'd10;
end

32'd322:
begin
    dest_x = `NOC_X_WIDTH'd2;
    dest_y = `NOC_Y_WIDTH'd10;
end

32'd323:
begin
    dest_x = `NOC_X_WIDTH'd3;
    dest_y = `NOC_Y_WIDTH'd10;
end

32'd324:
begin
    dest_x = `NOC_X_WIDTH'd4;
    dest_y = `NOC_Y_WIDTH'd10;
end

32'd325:
begin
    dest_x = `NOC_X_WIDTH'd5;
    dest_y = `NOC_Y_WIDTH'd10;
end

32'd326:
begin
    dest_x = `NOC_X_WIDTH'd6;
    dest_y = `NOC_Y_WIDTH'd10;
end

32'd327:
begin
    dest_x = `NOC_X_WIDTH'd7;
    dest_y = `NOC_Y_WIDTH'd10;
end

32'd328:
begin
    dest_x = `NOC_X_WIDTH'd8;
    dest_y = `NOC_Y_WIDTH'd10;
end

32'd329:
begin
    dest_x = `NOC_X_WIDTH'd9;
    dest_y = `NOC_Y_WIDTH'd10;
end

32'd330:
begin
    dest_x = `NOC_X_WIDTH'd10;
    dest_y = `NOC_Y_WIDTH'd10;
end

32'd331:
begin
    dest_x = `NOC_X_WIDTH'd11;
    dest_y = `NOC_Y_WIDTH'd10;
end

32'd332:
begin
    dest_x = `NOC_X_WIDTH'd12;
    dest_y = `NOC_Y_WIDTH'd10;
end

32'd333:
begin
    dest_x = `NOC_X_WIDTH'd13;
    dest_y = `NOC_Y_WIDTH'd10;
end

32'd334:
begin
    dest_x = `NOC_X_WIDTH'd14;
    dest_y = `NOC_Y_WIDTH'd10;
end

32'd335:
begin
    dest_x = `NOC_X_WIDTH'd15;
    dest_y = `NOC_Y_WIDTH'd10;
end

32'd336:
begin
    dest_x = `NOC_X_WIDTH'd16;
    dest_y = `NOC_Y_WIDTH'd10;
end

32'd337:
begin
    dest_x = `NOC_X_WIDTH'd17;
    dest_y = `NOC_Y_WIDTH'd10;
end

32'd338:
begin
    dest_x = `NOC_X_WIDTH'd18;
    dest_y = `NOC_Y_WIDTH'd10;
end

32'd339:
begin
    dest_x = `NOC_X_WIDTH'd19;
    dest_y = `NOC_Y_WIDTH'd10;
end

32'd340:
begin
    dest_x = `NOC_X_WIDTH'd20;
    dest_y = `NOC_Y_WIDTH'd10;
end

32'd341:
begin
    dest_x = `NOC_X_WIDTH'd21;
    dest_y = `NOC_Y_WIDTH'd10;
end

32'd342:
begin
    dest_x = `NOC_X_WIDTH'd22;
    dest_y = `NOC_Y_WIDTH'd10;
end

32'd343:
begin
    dest_x = `NOC_X_WIDTH'd23;
    dest_y = `NOC_Y_WIDTH'd10;
end

32'd344:
begin
    dest_x = `NOC_X_WIDTH'd24;
    dest_y = `NOC_Y_WIDTH'd10;
end

32'd345:
begin
    dest_x = `NOC_X_WIDTH'd25;
    dest_y = `NOC_Y_WIDTH'd10;
end

32'd346:
begin
    dest_x = `NOC_X_WIDTH'd26;
    dest_y = `NOC_Y_WIDTH'd10;
end

32'd347:
begin
    dest_x = `NOC_X_WIDTH'd27;
    dest_y = `NOC_Y_WIDTH'd10;
end

32'd348:
begin
    dest_x = `NOC_X_WIDTH'd28;
    dest_y = `NOC_Y_WIDTH'd10;
end

32'd349:
begin
    dest_x = `NOC_X_WIDTH'd29;
    dest_y = `NOC_Y_WIDTH'd10;
end

32'd350:
begin
    dest_x = `NOC_X_WIDTH'd30;
    dest_y = `NOC_Y_WIDTH'd10;
end

32'd351:
begin
    dest_x = `NOC_X_WIDTH'd31;
    dest_y = `NOC_Y_WIDTH'd10;
end

32'd352:
begin
    dest_x = `NOC_X_WIDTH'd0;
    dest_y = `NOC_Y_WIDTH'd11;
end

32'd353:
begin
    dest_x = `NOC_X_WIDTH'd1;
    dest_y = `NOC_Y_WIDTH'd11;
end

32'd354:
begin
    dest_x = `NOC_X_WIDTH'd2;
    dest_y = `NOC_Y_WIDTH'd11;
end

32'd355:
begin
    dest_x = `NOC_X_WIDTH'd3;
    dest_y = `NOC_Y_WIDTH'd11;
end

32'd356:
begin
    dest_x = `NOC_X_WIDTH'd4;
    dest_y = `NOC_Y_WIDTH'd11;
end

32'd357:
begin
    dest_x = `NOC_X_WIDTH'd5;
    dest_y = `NOC_Y_WIDTH'd11;
end

32'd358:
begin
    dest_x = `NOC_X_WIDTH'd6;
    dest_y = `NOC_Y_WIDTH'd11;
end

32'd359:
begin
    dest_x = `NOC_X_WIDTH'd7;
    dest_y = `NOC_Y_WIDTH'd11;
end

32'd360:
begin
    dest_x = `NOC_X_WIDTH'd8;
    dest_y = `NOC_Y_WIDTH'd11;
end

32'd361:
begin
    dest_x = `NOC_X_WIDTH'd9;
    dest_y = `NOC_Y_WIDTH'd11;
end

32'd362:
begin
    dest_x = `NOC_X_WIDTH'd10;
    dest_y = `NOC_Y_WIDTH'd11;
end

32'd363:
begin
    dest_x = `NOC_X_WIDTH'd11;
    dest_y = `NOC_Y_WIDTH'd11;
end

32'd364:
begin
    dest_x = `NOC_X_WIDTH'd12;
    dest_y = `NOC_Y_WIDTH'd11;
end

32'd365:
begin
    dest_x = `NOC_X_WIDTH'd13;
    dest_y = `NOC_Y_WIDTH'd11;
end

32'd366:
begin
    dest_x = `NOC_X_WIDTH'd14;
    dest_y = `NOC_Y_WIDTH'd11;
end

32'd367:
begin
    dest_x = `NOC_X_WIDTH'd15;
    dest_y = `NOC_Y_WIDTH'd11;
end

32'd368:
begin
    dest_x = `NOC_X_WIDTH'd16;
    dest_y = `NOC_Y_WIDTH'd11;
end

32'd369:
begin
    dest_x = `NOC_X_WIDTH'd17;
    dest_y = `NOC_Y_WIDTH'd11;
end

32'd370:
begin
    dest_x = `NOC_X_WIDTH'd18;
    dest_y = `NOC_Y_WIDTH'd11;
end

32'd371:
begin
    dest_x = `NOC_X_WIDTH'd19;
    dest_y = `NOC_Y_WIDTH'd11;
end

32'd372:
begin
    dest_x = `NOC_X_WIDTH'd20;
    dest_y = `NOC_Y_WIDTH'd11;
end

32'd373:
begin
    dest_x = `NOC_X_WIDTH'd21;
    dest_y = `NOC_Y_WIDTH'd11;
end

32'd374:
begin
    dest_x = `NOC_X_WIDTH'd22;
    dest_y = `NOC_Y_WIDTH'd11;
end

32'd375:
begin
    dest_x = `NOC_X_WIDTH'd23;
    dest_y = `NOC_Y_WIDTH'd11;
end

32'd376:
begin
    dest_x = `NOC_X_WIDTH'd24;
    dest_y = `NOC_Y_WIDTH'd11;
end

32'd377:
begin
    dest_x = `NOC_X_WIDTH'd25;
    dest_y = `NOC_Y_WIDTH'd11;
end

32'd378:
begin
    dest_x = `NOC_X_WIDTH'd26;
    dest_y = `NOC_Y_WIDTH'd11;
end

32'd379:
begin
    dest_x = `NOC_X_WIDTH'd27;
    dest_y = `NOC_Y_WIDTH'd11;
end

32'd380:
begin
    dest_x = `NOC_X_WIDTH'd28;
    dest_y = `NOC_Y_WIDTH'd11;
end

32'd381:
begin
    dest_x = `NOC_X_WIDTH'd29;
    dest_y = `NOC_Y_WIDTH'd11;
end

32'd382:
begin
    dest_x = `NOC_X_WIDTH'd30;
    dest_y = `NOC_Y_WIDTH'd11;
end

32'd383:
begin
    dest_x = `NOC_X_WIDTH'd31;
    dest_y = `NOC_Y_WIDTH'd11;
end

32'd384:
begin
    dest_x = `NOC_X_WIDTH'd0;
    dest_y = `NOC_Y_WIDTH'd12;
end

32'd385:
begin
    dest_x = `NOC_X_WIDTH'd1;
    dest_y = `NOC_Y_WIDTH'd12;
end

32'd386:
begin
    dest_x = `NOC_X_WIDTH'd2;
    dest_y = `NOC_Y_WIDTH'd12;
end

32'd387:
begin
    dest_x = `NOC_X_WIDTH'd3;
    dest_y = `NOC_Y_WIDTH'd12;
end

32'd388:
begin
    dest_x = `NOC_X_WIDTH'd4;
    dest_y = `NOC_Y_WIDTH'd12;
end

32'd389:
begin
    dest_x = `NOC_X_WIDTH'd5;
    dest_y = `NOC_Y_WIDTH'd12;
end

32'd390:
begin
    dest_x = `NOC_X_WIDTH'd6;
    dest_y = `NOC_Y_WIDTH'd12;
end

32'd391:
begin
    dest_x = `NOC_X_WIDTH'd7;
    dest_y = `NOC_Y_WIDTH'd12;
end

32'd392:
begin
    dest_x = `NOC_X_WIDTH'd8;
    dest_y = `NOC_Y_WIDTH'd12;
end

32'd393:
begin
    dest_x = `NOC_X_WIDTH'd9;
    dest_y = `NOC_Y_WIDTH'd12;
end

32'd394:
begin
    dest_x = `NOC_X_WIDTH'd10;
    dest_y = `NOC_Y_WIDTH'd12;
end

32'd395:
begin
    dest_x = `NOC_X_WIDTH'd11;
    dest_y = `NOC_Y_WIDTH'd12;
end

32'd396:
begin
    dest_x = `NOC_X_WIDTH'd12;
    dest_y = `NOC_Y_WIDTH'd12;
end

32'd397:
begin
    dest_x = `NOC_X_WIDTH'd13;
    dest_y = `NOC_Y_WIDTH'd12;
end

32'd398:
begin
    dest_x = `NOC_X_WIDTH'd14;
    dest_y = `NOC_Y_WIDTH'd12;
end

32'd399:
begin
    dest_x = `NOC_X_WIDTH'd15;
    dest_y = `NOC_Y_WIDTH'd12;
end

32'd400:
begin
    dest_x = `NOC_X_WIDTH'd16;
    dest_y = `NOC_Y_WIDTH'd12;
end

32'd401:
begin
    dest_x = `NOC_X_WIDTH'd17;
    dest_y = `NOC_Y_WIDTH'd12;
end

32'd402:
begin
    dest_x = `NOC_X_WIDTH'd18;
    dest_y = `NOC_Y_WIDTH'd12;
end

32'd403:
begin
    dest_x = `NOC_X_WIDTH'd19;
    dest_y = `NOC_Y_WIDTH'd12;
end

32'd404:
begin
    dest_x = `NOC_X_WIDTH'd20;
    dest_y = `NOC_Y_WIDTH'd12;
end

32'd405:
begin
    dest_x = `NOC_X_WIDTH'd21;
    dest_y = `NOC_Y_WIDTH'd12;
end

32'd406:
begin
    dest_x = `NOC_X_WIDTH'd22;
    dest_y = `NOC_Y_WIDTH'd12;
end

32'd407:
begin
    dest_x = `NOC_X_WIDTH'd23;
    dest_y = `NOC_Y_WIDTH'd12;
end

32'd408:
begin
    dest_x = `NOC_X_WIDTH'd24;
    dest_y = `NOC_Y_WIDTH'd12;
end

32'd409:
begin
    dest_x = `NOC_X_WIDTH'd25;
    dest_y = `NOC_Y_WIDTH'd12;
end

32'd410:
begin
    dest_x = `NOC_X_WIDTH'd26;
    dest_y = `NOC_Y_WIDTH'd12;
end

32'd411:
begin
    dest_x = `NOC_X_WIDTH'd27;
    dest_y = `NOC_Y_WIDTH'd12;
end

32'd412:
begin
    dest_x = `NOC_X_WIDTH'd28;
    dest_y = `NOC_Y_WIDTH'd12;
end

32'd413:
begin
    dest_x = `NOC_X_WIDTH'd29;
    dest_y = `NOC_Y_WIDTH'd12;
end

32'd414:
begin
    dest_x = `NOC_X_WIDTH'd30;
    dest_y = `NOC_Y_WIDTH'd12;
end

32'd415:
begin
    dest_x = `NOC_X_WIDTH'd31;
    dest_y = `NOC_Y_WIDTH'd12;
end

32'd416:
begin
    dest_x = `NOC_X_WIDTH'd0;
    dest_y = `NOC_Y_WIDTH'd13;
end

32'd417:
begin
    dest_x = `NOC_X_WIDTH'd1;
    dest_y = `NOC_Y_WIDTH'd13;
end

32'd418:
begin
    dest_x = `NOC_X_WIDTH'd2;
    dest_y = `NOC_Y_WIDTH'd13;
end

32'd419:
begin
    dest_x = `NOC_X_WIDTH'd3;
    dest_y = `NOC_Y_WIDTH'd13;
end

32'd420:
begin
    dest_x = `NOC_X_WIDTH'd4;
    dest_y = `NOC_Y_WIDTH'd13;
end

32'd421:
begin
    dest_x = `NOC_X_WIDTH'd5;
    dest_y = `NOC_Y_WIDTH'd13;
end

32'd422:
begin
    dest_x = `NOC_X_WIDTH'd6;
    dest_y = `NOC_Y_WIDTH'd13;
end

32'd423:
begin
    dest_x = `NOC_X_WIDTH'd7;
    dest_y = `NOC_Y_WIDTH'd13;
end

32'd424:
begin
    dest_x = `NOC_X_WIDTH'd8;
    dest_y = `NOC_Y_WIDTH'd13;
end

32'd425:
begin
    dest_x = `NOC_X_WIDTH'd9;
    dest_y = `NOC_Y_WIDTH'd13;
end

32'd426:
begin
    dest_x = `NOC_X_WIDTH'd10;
    dest_y = `NOC_Y_WIDTH'd13;
end

32'd427:
begin
    dest_x = `NOC_X_WIDTH'd11;
    dest_y = `NOC_Y_WIDTH'd13;
end

32'd428:
begin
    dest_x = `NOC_X_WIDTH'd12;
    dest_y = `NOC_Y_WIDTH'd13;
end

32'd429:
begin
    dest_x = `NOC_X_WIDTH'd13;
    dest_y = `NOC_Y_WIDTH'd13;
end

32'd430:
begin
    dest_x = `NOC_X_WIDTH'd14;
    dest_y = `NOC_Y_WIDTH'd13;
end

32'd431:
begin
    dest_x = `NOC_X_WIDTH'd15;
    dest_y = `NOC_Y_WIDTH'd13;
end

32'd432:
begin
    dest_x = `NOC_X_WIDTH'd16;
    dest_y = `NOC_Y_WIDTH'd13;
end

32'd433:
begin
    dest_x = `NOC_X_WIDTH'd17;
    dest_y = `NOC_Y_WIDTH'd13;
end

32'd434:
begin
    dest_x = `NOC_X_WIDTH'd18;
    dest_y = `NOC_Y_WIDTH'd13;
end

32'd435:
begin
    dest_x = `NOC_X_WIDTH'd19;
    dest_y = `NOC_Y_WIDTH'd13;
end

32'd436:
begin
    dest_x = `NOC_X_WIDTH'd20;
    dest_y = `NOC_Y_WIDTH'd13;
end

32'd437:
begin
    dest_x = `NOC_X_WIDTH'd21;
    dest_y = `NOC_Y_WIDTH'd13;
end

32'd438:
begin
    dest_x = `NOC_X_WIDTH'd22;
    dest_y = `NOC_Y_WIDTH'd13;
end

32'd439:
begin
    dest_x = `NOC_X_WIDTH'd23;
    dest_y = `NOC_Y_WIDTH'd13;
end

32'd440:
begin
    dest_x = `NOC_X_WIDTH'd24;
    dest_y = `NOC_Y_WIDTH'd13;
end

32'd441:
begin
    dest_x = `NOC_X_WIDTH'd25;
    dest_y = `NOC_Y_WIDTH'd13;
end

32'd442:
begin
    dest_x = `NOC_X_WIDTH'd26;
    dest_y = `NOC_Y_WIDTH'd13;
end

32'd443:
begin
    dest_x = `NOC_X_WIDTH'd27;
    dest_y = `NOC_Y_WIDTH'd13;
end

32'd444:
begin
    dest_x = `NOC_X_WIDTH'd28;
    dest_y = `NOC_Y_WIDTH'd13;
end

32'd445:
begin
    dest_x = `NOC_X_WIDTH'd29;
    dest_y = `NOC_Y_WIDTH'd13;
end

32'd446:
begin
    dest_x = `NOC_X_WIDTH'd30;
    dest_y = `NOC_Y_WIDTH'd13;
end

32'd447:
begin
    dest_x = `NOC_X_WIDTH'd31;
    dest_y = `NOC_Y_WIDTH'd13;
end

32'd448:
begin
    dest_x = `NOC_X_WIDTH'd0;
    dest_y = `NOC_Y_WIDTH'd14;
end

32'd449:
begin
    dest_x = `NOC_X_WIDTH'd1;
    dest_y = `NOC_Y_WIDTH'd14;
end

32'd450:
begin
    dest_x = `NOC_X_WIDTH'd2;
    dest_y = `NOC_Y_WIDTH'd14;
end

32'd451:
begin
    dest_x = `NOC_X_WIDTH'd3;
    dest_y = `NOC_Y_WIDTH'd14;
end

32'd452:
begin
    dest_x = `NOC_X_WIDTH'd4;
    dest_y = `NOC_Y_WIDTH'd14;
end

32'd453:
begin
    dest_x = `NOC_X_WIDTH'd5;
    dest_y = `NOC_Y_WIDTH'd14;
end

32'd454:
begin
    dest_x = `NOC_X_WIDTH'd6;
    dest_y = `NOC_Y_WIDTH'd14;
end

32'd455:
begin
    dest_x = `NOC_X_WIDTH'd7;
    dest_y = `NOC_Y_WIDTH'd14;
end

32'd456:
begin
    dest_x = `NOC_X_WIDTH'd8;
    dest_y = `NOC_Y_WIDTH'd14;
end

32'd457:
begin
    dest_x = `NOC_X_WIDTH'd9;
    dest_y = `NOC_Y_WIDTH'd14;
end

32'd458:
begin
    dest_x = `NOC_X_WIDTH'd10;
    dest_y = `NOC_Y_WIDTH'd14;
end

32'd459:
begin
    dest_x = `NOC_X_WIDTH'd11;
    dest_y = `NOC_Y_WIDTH'd14;
end

32'd460:
begin
    dest_x = `NOC_X_WIDTH'd12;
    dest_y = `NOC_Y_WIDTH'd14;
end

32'd461:
begin
    dest_x = `NOC_X_WIDTH'd13;
    dest_y = `NOC_Y_WIDTH'd14;
end

32'd462:
begin
    dest_x = `NOC_X_WIDTH'd14;
    dest_y = `NOC_Y_WIDTH'd14;
end

32'd463:
begin
    dest_x = `NOC_X_WIDTH'd15;
    dest_y = `NOC_Y_WIDTH'd14;
end

32'd464:
begin
    dest_x = `NOC_X_WIDTH'd16;
    dest_y = `NOC_Y_WIDTH'd14;
end

32'd465:
begin
    dest_x = `NOC_X_WIDTH'd17;
    dest_y = `NOC_Y_WIDTH'd14;
end

32'd466:
begin
    dest_x = `NOC_X_WIDTH'd18;
    dest_y = `NOC_Y_WIDTH'd14;
end

32'd467:
begin
    dest_x = `NOC_X_WIDTH'd19;
    dest_y = `NOC_Y_WIDTH'd14;
end

32'd468:
begin
    dest_x = `NOC_X_WIDTH'd20;
    dest_y = `NOC_Y_WIDTH'd14;
end

32'd469:
begin
    dest_x = `NOC_X_WIDTH'd21;
    dest_y = `NOC_Y_WIDTH'd14;
end

32'd470:
begin
    dest_x = `NOC_X_WIDTH'd22;
    dest_y = `NOC_Y_WIDTH'd14;
end

32'd471:
begin
    dest_x = `NOC_X_WIDTH'd23;
    dest_y = `NOC_Y_WIDTH'd14;
end

32'd472:
begin
    dest_x = `NOC_X_WIDTH'd24;
    dest_y = `NOC_Y_WIDTH'd14;
end

32'd473:
begin
    dest_x = `NOC_X_WIDTH'd25;
    dest_y = `NOC_Y_WIDTH'd14;
end

32'd474:
begin
    dest_x = `NOC_X_WIDTH'd26;
    dest_y = `NOC_Y_WIDTH'd14;
end

32'd475:
begin
    dest_x = `NOC_X_WIDTH'd27;
    dest_y = `NOC_Y_WIDTH'd14;
end

32'd476:
begin
    dest_x = `NOC_X_WIDTH'd28;
    dest_y = `NOC_Y_WIDTH'd14;
end

32'd477:
begin
    dest_x = `NOC_X_WIDTH'd29;
    dest_y = `NOC_Y_WIDTH'd14;
end

32'd478:
begin
    dest_x = `NOC_X_WIDTH'd30;
    dest_y = `NOC_Y_WIDTH'd14;
end

32'd479:
begin
    dest_x = `NOC_X_WIDTH'd31;
    dest_y = `NOC_Y_WIDTH'd14;
end

32'd480:
begin
    dest_x = `NOC_X_WIDTH'd0;
    dest_y = `NOC_Y_WIDTH'd15;
end

32'd481:
begin
    dest_x = `NOC_X_WIDTH'd1;
    dest_y = `NOC_Y_WIDTH'd15;
end

32'd482:
begin
    dest_x = `NOC_X_WIDTH'd2;
    dest_y = `NOC_Y_WIDTH'd15;
end

32'd483:
begin
    dest_x = `NOC_X_WIDTH'd3;
    dest_y = `NOC_Y_WIDTH'd15;
end

32'd484:
begin
    dest_x = `NOC_X_WIDTH'd4;
    dest_y = `NOC_Y_WIDTH'd15;
end

32'd485:
begin
    dest_x = `NOC_X_WIDTH'd5;
    dest_y = `NOC_Y_WIDTH'd15;
end

32'd486:
begin
    dest_x = `NOC_X_WIDTH'd6;
    dest_y = `NOC_Y_WIDTH'd15;
end

32'd487:
begin
    dest_x = `NOC_X_WIDTH'd7;
    dest_y = `NOC_Y_WIDTH'd15;
end

32'd488:
begin
    dest_x = `NOC_X_WIDTH'd8;
    dest_y = `NOC_Y_WIDTH'd15;
end

32'd489:
begin
    dest_x = `NOC_X_WIDTH'd9;
    dest_y = `NOC_Y_WIDTH'd15;
end

32'd490:
begin
    dest_x = `NOC_X_WIDTH'd10;
    dest_y = `NOC_Y_WIDTH'd15;
end

32'd491:
begin
    dest_x = `NOC_X_WIDTH'd11;
    dest_y = `NOC_Y_WIDTH'd15;
end

32'd492:
begin
    dest_x = `NOC_X_WIDTH'd12;
    dest_y = `NOC_Y_WIDTH'd15;
end

32'd493:
begin
    dest_x = `NOC_X_WIDTH'd13;
    dest_y = `NOC_Y_WIDTH'd15;
end

32'd494:
begin
    dest_x = `NOC_X_WIDTH'd14;
    dest_y = `NOC_Y_WIDTH'd15;
end

32'd495:
begin
    dest_x = `NOC_X_WIDTH'd15;
    dest_y = `NOC_Y_WIDTH'd15;
end

32'd496:
begin
    dest_x = `NOC_X_WIDTH'd16;
    dest_y = `NOC_Y_WIDTH'd15;
end

32'd497:
begin
    dest_x = `NOC_X_WIDTH'd17;
    dest_y = `NOC_Y_WIDTH'd15;
end

32'd498:
begin
    dest_x = `NOC_X_WIDTH'd18;
    dest_y = `NOC_Y_WIDTH'd15;
end

32'd499:
begin
    dest_x = `NOC_X_WIDTH'd19;
    dest_y = `NOC_Y_WIDTH'd15;
end

32'd500:
begin
    dest_x = `NOC_X_WIDTH'd20;
    dest_y = `NOC_Y_WIDTH'd15;
end

32'd501:
begin
    dest_x = `NOC_X_WIDTH'd21;
    dest_y = `NOC_Y_WIDTH'd15;
end

32'd502:
begin
    dest_x = `NOC_X_WIDTH'd22;
    dest_y = `NOC_Y_WIDTH'd15;
end

32'd503:
begin
    dest_x = `NOC_X_WIDTH'd23;
    dest_y = `NOC_Y_WIDTH'd15;
end

32'd504:
begin
    dest_x = `NOC_X_WIDTH'd24;
    dest_y = `NOC_Y_WIDTH'd15;
end

32'd505:
begin
    dest_x = `NOC_X_WIDTH'd25;
    dest_y = `NOC_Y_WIDTH'd15;
end

32'd506:
begin
    dest_x = `NOC_X_WIDTH'd26;
    dest_y = `NOC_Y_WIDTH'd15;
end

32'd507:
begin
    dest_x = `NOC_X_WIDTH'd27;
    dest_y = `NOC_Y_WIDTH'd15;
end

32'd508:
begin
    dest_x = `NOC_X_WIDTH'd28;
    dest_y = `NOC_Y_WIDTH'd15;
end

32'd509:
begin
    dest_x = `NOC_X_WIDTH'd29;
    dest_y = `NOC_Y_WIDTH'd15;
end

32'd510:
begin
    dest_x = `NOC_X_WIDTH'd30;
    dest_y = `NOC_Y_WIDTH'd15;
end

32'd511:
begin
    dest_x = `NOC_X_WIDTH'd31;
    dest_y = `NOC_Y_WIDTH'd15;
end

32'd512:
begin
    dest_x = `NOC_X_WIDTH'd0;
    dest_y = `NOC_Y_WIDTH'd16;
end

32'd513:
begin
    dest_x = `NOC_X_WIDTH'd1;
    dest_y = `NOC_Y_WIDTH'd16;
end

32'd514:
begin
    dest_x = `NOC_X_WIDTH'd2;
    dest_y = `NOC_Y_WIDTH'd16;
end

32'd515:
begin
    dest_x = `NOC_X_WIDTH'd3;
    dest_y = `NOC_Y_WIDTH'd16;
end

32'd516:
begin
    dest_x = `NOC_X_WIDTH'd4;
    dest_y = `NOC_Y_WIDTH'd16;
end

32'd517:
begin
    dest_x = `NOC_X_WIDTH'd5;
    dest_y = `NOC_Y_WIDTH'd16;
end

32'd518:
begin
    dest_x = `NOC_X_WIDTH'd6;
    dest_y = `NOC_Y_WIDTH'd16;
end

32'd519:
begin
    dest_x = `NOC_X_WIDTH'd7;
    dest_y = `NOC_Y_WIDTH'd16;
end

32'd520:
begin
    dest_x = `NOC_X_WIDTH'd8;
    dest_y = `NOC_Y_WIDTH'd16;
end

32'd521:
begin
    dest_x = `NOC_X_WIDTH'd9;
    dest_y = `NOC_Y_WIDTH'd16;
end

32'd522:
begin
    dest_x = `NOC_X_WIDTH'd10;
    dest_y = `NOC_Y_WIDTH'd16;
end

32'd523:
begin
    dest_x = `NOC_X_WIDTH'd11;
    dest_y = `NOC_Y_WIDTH'd16;
end

32'd524:
begin
    dest_x = `NOC_X_WIDTH'd12;
    dest_y = `NOC_Y_WIDTH'd16;
end

32'd525:
begin
    dest_x = `NOC_X_WIDTH'd13;
    dest_y = `NOC_Y_WIDTH'd16;
end

32'd526:
begin
    dest_x = `NOC_X_WIDTH'd14;
    dest_y = `NOC_Y_WIDTH'd16;
end

32'd527:
begin
    dest_x = `NOC_X_WIDTH'd15;
    dest_y = `NOC_Y_WIDTH'd16;
end

32'd528:
begin
    dest_x = `NOC_X_WIDTH'd16;
    dest_y = `NOC_Y_WIDTH'd16;
end

32'd529:
begin
    dest_x = `NOC_X_WIDTH'd17;
    dest_y = `NOC_Y_WIDTH'd16;
end

32'd530:
begin
    dest_x = `NOC_X_WIDTH'd18;
    dest_y = `NOC_Y_WIDTH'd16;
end

32'd531:
begin
    dest_x = `NOC_X_WIDTH'd19;
    dest_y = `NOC_Y_WIDTH'd16;
end

32'd532:
begin
    dest_x = `NOC_X_WIDTH'd20;
    dest_y = `NOC_Y_WIDTH'd16;
end

32'd533:
begin
    dest_x = `NOC_X_WIDTH'd21;
    dest_y = `NOC_Y_WIDTH'd16;
end

32'd534:
begin
    dest_x = `NOC_X_WIDTH'd22;
    dest_y = `NOC_Y_WIDTH'd16;
end

32'd535:
begin
    dest_x = `NOC_X_WIDTH'd23;
    dest_y = `NOC_Y_WIDTH'd16;
end

32'd536:
begin
    dest_x = `NOC_X_WIDTH'd24;
    dest_y = `NOC_Y_WIDTH'd16;
end

32'd537:
begin
    dest_x = `NOC_X_WIDTH'd25;
    dest_y = `NOC_Y_WIDTH'd16;
end

32'd538:
begin
    dest_x = `NOC_X_WIDTH'd26;
    dest_y = `NOC_Y_WIDTH'd16;
end

32'd539:
begin
    dest_x = `NOC_X_WIDTH'd27;
    dest_y = `NOC_Y_WIDTH'd16;
end

32'd540:
begin
    dest_x = `NOC_X_WIDTH'd28;
    dest_y = `NOC_Y_WIDTH'd16;
end

32'd541:
begin
    dest_x = `NOC_X_WIDTH'd29;
    dest_y = `NOC_Y_WIDTH'd16;
end

32'd542:
begin
    dest_x = `NOC_X_WIDTH'd30;
    dest_y = `NOC_Y_WIDTH'd16;
end

32'd543:
begin
    dest_x = `NOC_X_WIDTH'd31;
    dest_y = `NOC_Y_WIDTH'd16;
end

32'd544:
begin
    dest_x = `NOC_X_WIDTH'd0;
    dest_y = `NOC_Y_WIDTH'd17;
end

32'd545:
begin
    dest_x = `NOC_X_WIDTH'd1;
    dest_y = `NOC_Y_WIDTH'd17;
end

32'd546:
begin
    dest_x = `NOC_X_WIDTH'd2;
    dest_y = `NOC_Y_WIDTH'd17;
end

32'd547:
begin
    dest_x = `NOC_X_WIDTH'd3;
    dest_y = `NOC_Y_WIDTH'd17;
end

32'd548:
begin
    dest_x = `NOC_X_WIDTH'd4;
    dest_y = `NOC_Y_WIDTH'd17;
end

32'd549:
begin
    dest_x = `NOC_X_WIDTH'd5;
    dest_y = `NOC_Y_WIDTH'd17;
end

32'd550:
begin
    dest_x = `NOC_X_WIDTH'd6;
    dest_y = `NOC_Y_WIDTH'd17;
end

32'd551:
begin
    dest_x = `NOC_X_WIDTH'd7;
    dest_y = `NOC_Y_WIDTH'd17;
end

32'd552:
begin
    dest_x = `NOC_X_WIDTH'd8;
    dest_y = `NOC_Y_WIDTH'd17;
end

32'd553:
begin
    dest_x = `NOC_X_WIDTH'd9;
    dest_y = `NOC_Y_WIDTH'd17;
end

32'd554:
begin
    dest_x = `NOC_X_WIDTH'd10;
    dest_y = `NOC_Y_WIDTH'd17;
end

32'd555:
begin
    dest_x = `NOC_X_WIDTH'd11;
    dest_y = `NOC_Y_WIDTH'd17;
end

32'd556:
begin
    dest_x = `NOC_X_WIDTH'd12;
    dest_y = `NOC_Y_WIDTH'd17;
end

32'd557:
begin
    dest_x = `NOC_X_WIDTH'd13;
    dest_y = `NOC_Y_WIDTH'd17;
end

32'd558:
begin
    dest_x = `NOC_X_WIDTH'd14;
    dest_y = `NOC_Y_WIDTH'd17;
end

32'd559:
begin
    dest_x = `NOC_X_WIDTH'd15;
    dest_y = `NOC_Y_WIDTH'd17;
end

32'd560:
begin
    dest_x = `NOC_X_WIDTH'd16;
    dest_y = `NOC_Y_WIDTH'd17;
end

32'd561:
begin
    dest_x = `NOC_X_WIDTH'd17;
    dest_y = `NOC_Y_WIDTH'd17;
end

32'd562:
begin
    dest_x = `NOC_X_WIDTH'd18;
    dest_y = `NOC_Y_WIDTH'd17;
end

32'd563:
begin
    dest_x = `NOC_X_WIDTH'd19;
    dest_y = `NOC_Y_WIDTH'd17;
end

32'd564:
begin
    dest_x = `NOC_X_WIDTH'd20;
    dest_y = `NOC_Y_WIDTH'd17;
end

32'd565:
begin
    dest_x = `NOC_X_WIDTH'd21;
    dest_y = `NOC_Y_WIDTH'd17;
end

32'd566:
begin
    dest_x = `NOC_X_WIDTH'd22;
    dest_y = `NOC_Y_WIDTH'd17;
end

32'd567:
begin
    dest_x = `NOC_X_WIDTH'd23;
    dest_y = `NOC_Y_WIDTH'd17;
end

32'd568:
begin
    dest_x = `NOC_X_WIDTH'd24;
    dest_y = `NOC_Y_WIDTH'd17;
end

32'd569:
begin
    dest_x = `NOC_X_WIDTH'd25;
    dest_y = `NOC_Y_WIDTH'd17;
end

32'd570:
begin
    dest_x = `NOC_X_WIDTH'd26;
    dest_y = `NOC_Y_WIDTH'd17;
end

32'd571:
begin
    dest_x = `NOC_X_WIDTH'd27;
    dest_y = `NOC_Y_WIDTH'd17;
end

32'd572:
begin
    dest_x = `NOC_X_WIDTH'd28;
    dest_y = `NOC_Y_WIDTH'd17;
end

32'd573:
begin
    dest_x = `NOC_X_WIDTH'd29;
    dest_y = `NOC_Y_WIDTH'd17;
end

32'd574:
begin
    dest_x = `NOC_X_WIDTH'd30;
    dest_y = `NOC_Y_WIDTH'd17;
end

32'd575:
begin
    dest_x = `NOC_X_WIDTH'd31;
    dest_y = `NOC_Y_WIDTH'd17;
end

32'd576:
begin
    dest_x = `NOC_X_WIDTH'd0;
    dest_y = `NOC_Y_WIDTH'd18;
end

32'd577:
begin
    dest_x = `NOC_X_WIDTH'd1;
    dest_y = `NOC_Y_WIDTH'd18;
end

32'd578:
begin
    dest_x = `NOC_X_WIDTH'd2;
    dest_y = `NOC_Y_WIDTH'd18;
end

32'd579:
begin
    dest_x = `NOC_X_WIDTH'd3;
    dest_y = `NOC_Y_WIDTH'd18;
end

32'd580:
begin
    dest_x = `NOC_X_WIDTH'd4;
    dest_y = `NOC_Y_WIDTH'd18;
end

32'd581:
begin
    dest_x = `NOC_X_WIDTH'd5;
    dest_y = `NOC_Y_WIDTH'd18;
end

32'd582:
begin
    dest_x = `NOC_X_WIDTH'd6;
    dest_y = `NOC_Y_WIDTH'd18;
end

32'd583:
begin
    dest_x = `NOC_X_WIDTH'd7;
    dest_y = `NOC_Y_WIDTH'd18;
end

32'd584:
begin
    dest_x = `NOC_X_WIDTH'd8;
    dest_y = `NOC_Y_WIDTH'd18;
end

32'd585:
begin
    dest_x = `NOC_X_WIDTH'd9;
    dest_y = `NOC_Y_WIDTH'd18;
end

32'd586:
begin
    dest_x = `NOC_X_WIDTH'd10;
    dest_y = `NOC_Y_WIDTH'd18;
end

32'd587:
begin
    dest_x = `NOC_X_WIDTH'd11;
    dest_y = `NOC_Y_WIDTH'd18;
end

32'd588:
begin
    dest_x = `NOC_X_WIDTH'd12;
    dest_y = `NOC_Y_WIDTH'd18;
end

32'd589:
begin
    dest_x = `NOC_X_WIDTH'd13;
    dest_y = `NOC_Y_WIDTH'd18;
end

32'd590:
begin
    dest_x = `NOC_X_WIDTH'd14;
    dest_y = `NOC_Y_WIDTH'd18;
end

32'd591:
begin
    dest_x = `NOC_X_WIDTH'd15;
    dest_y = `NOC_Y_WIDTH'd18;
end

32'd592:
begin
    dest_x = `NOC_X_WIDTH'd16;
    dest_y = `NOC_Y_WIDTH'd18;
end

32'd593:
begin
    dest_x = `NOC_X_WIDTH'd17;
    dest_y = `NOC_Y_WIDTH'd18;
end

32'd594:
begin
    dest_x = `NOC_X_WIDTH'd18;
    dest_y = `NOC_Y_WIDTH'd18;
end

32'd595:
begin
    dest_x = `NOC_X_WIDTH'd19;
    dest_y = `NOC_Y_WIDTH'd18;
end

32'd596:
begin
    dest_x = `NOC_X_WIDTH'd20;
    dest_y = `NOC_Y_WIDTH'd18;
end

32'd597:
begin
    dest_x = `NOC_X_WIDTH'd21;
    dest_y = `NOC_Y_WIDTH'd18;
end

32'd598:
begin
    dest_x = `NOC_X_WIDTH'd22;
    dest_y = `NOC_Y_WIDTH'd18;
end

32'd599:
begin
    dest_x = `NOC_X_WIDTH'd23;
    dest_y = `NOC_Y_WIDTH'd18;
end

32'd600:
begin
    dest_x = `NOC_X_WIDTH'd24;
    dest_y = `NOC_Y_WIDTH'd18;
end

32'd601:
begin
    dest_x = `NOC_X_WIDTH'd25;
    dest_y = `NOC_Y_WIDTH'd18;
end

32'd602:
begin
    dest_x = `NOC_X_WIDTH'd26;
    dest_y = `NOC_Y_WIDTH'd18;
end

32'd603:
begin
    dest_x = `NOC_X_WIDTH'd27;
    dest_y = `NOC_Y_WIDTH'd18;
end

32'd604:
begin
    dest_x = `NOC_X_WIDTH'd28;
    dest_y = `NOC_Y_WIDTH'd18;
end

32'd605:
begin
    dest_x = `NOC_X_WIDTH'd29;
    dest_y = `NOC_Y_WIDTH'd18;
end

32'd606:
begin
    dest_x = `NOC_X_WIDTH'd30;
    dest_y = `NOC_Y_WIDTH'd18;
end

32'd607:
begin
    dest_x = `NOC_X_WIDTH'd31;
    dest_y = `NOC_Y_WIDTH'd18;
end

32'd608:
begin
    dest_x = `NOC_X_WIDTH'd0;
    dest_y = `NOC_Y_WIDTH'd19;
end

32'd609:
begin
    dest_x = `NOC_X_WIDTH'd1;
    dest_y = `NOC_Y_WIDTH'd19;
end

32'd610:
begin
    dest_x = `NOC_X_WIDTH'd2;
    dest_y = `NOC_Y_WIDTH'd19;
end

32'd611:
begin
    dest_x = `NOC_X_WIDTH'd3;
    dest_y = `NOC_Y_WIDTH'd19;
end

32'd612:
begin
    dest_x = `NOC_X_WIDTH'd4;
    dest_y = `NOC_Y_WIDTH'd19;
end

32'd613:
begin
    dest_x = `NOC_X_WIDTH'd5;
    dest_y = `NOC_Y_WIDTH'd19;
end

32'd614:
begin
    dest_x = `NOC_X_WIDTH'd6;
    dest_y = `NOC_Y_WIDTH'd19;
end

32'd615:
begin
    dest_x = `NOC_X_WIDTH'd7;
    dest_y = `NOC_Y_WIDTH'd19;
end

32'd616:
begin
    dest_x = `NOC_X_WIDTH'd8;
    dest_y = `NOC_Y_WIDTH'd19;
end

32'd617:
begin
    dest_x = `NOC_X_WIDTH'd9;
    dest_y = `NOC_Y_WIDTH'd19;
end

32'd618:
begin
    dest_x = `NOC_X_WIDTH'd10;
    dest_y = `NOC_Y_WIDTH'd19;
end

32'd619:
begin
    dest_x = `NOC_X_WIDTH'd11;
    dest_y = `NOC_Y_WIDTH'd19;
end

32'd620:
begin
    dest_x = `NOC_X_WIDTH'd12;
    dest_y = `NOC_Y_WIDTH'd19;
end

32'd621:
begin
    dest_x = `NOC_X_WIDTH'd13;
    dest_y = `NOC_Y_WIDTH'd19;
end

32'd622:
begin
    dest_x = `NOC_X_WIDTH'd14;
    dest_y = `NOC_Y_WIDTH'd19;
end

32'd623:
begin
    dest_x = `NOC_X_WIDTH'd15;
    dest_y = `NOC_Y_WIDTH'd19;
end

32'd624:
begin
    dest_x = `NOC_X_WIDTH'd16;
    dest_y = `NOC_Y_WIDTH'd19;
end

32'd625:
begin
    dest_x = `NOC_X_WIDTH'd17;
    dest_y = `NOC_Y_WIDTH'd19;
end

32'd626:
begin
    dest_x = `NOC_X_WIDTH'd18;
    dest_y = `NOC_Y_WIDTH'd19;
end

32'd627:
begin
    dest_x = `NOC_X_WIDTH'd19;
    dest_y = `NOC_Y_WIDTH'd19;
end

32'd628:
begin
    dest_x = `NOC_X_WIDTH'd20;
    dest_y = `NOC_Y_WIDTH'd19;
end

32'd629:
begin
    dest_x = `NOC_X_WIDTH'd21;
    dest_y = `NOC_Y_WIDTH'd19;
end

32'd630:
begin
    dest_x = `NOC_X_WIDTH'd22;
    dest_y = `NOC_Y_WIDTH'd19;
end

32'd631:
begin
    dest_x = `NOC_X_WIDTH'd23;
    dest_y = `NOC_Y_WIDTH'd19;
end

32'd632:
begin
    dest_x = `NOC_X_WIDTH'd24;
    dest_y = `NOC_Y_WIDTH'd19;
end

32'd633:
begin
    dest_x = `NOC_X_WIDTH'd25;
    dest_y = `NOC_Y_WIDTH'd19;
end

32'd634:
begin
    dest_x = `NOC_X_WIDTH'd26;
    dest_y = `NOC_Y_WIDTH'd19;
end

32'd635:
begin
    dest_x = `NOC_X_WIDTH'd27;
    dest_y = `NOC_Y_WIDTH'd19;
end

32'd636:
begin
    dest_x = `NOC_X_WIDTH'd28;
    dest_y = `NOC_Y_WIDTH'd19;
end

32'd637:
begin
    dest_x = `NOC_X_WIDTH'd29;
    dest_y = `NOC_Y_WIDTH'd19;
end

32'd638:
begin
    dest_x = `NOC_X_WIDTH'd30;
    dest_y = `NOC_Y_WIDTH'd19;
end

32'd639:
begin
    dest_x = `NOC_X_WIDTH'd31;
    dest_y = `NOC_Y_WIDTH'd19;
end

32'd640:
begin
    dest_x = `NOC_X_WIDTH'd0;
    dest_y = `NOC_Y_WIDTH'd20;
end

32'd641:
begin
    dest_x = `NOC_X_WIDTH'd1;
    dest_y = `NOC_Y_WIDTH'd20;
end

32'd642:
begin
    dest_x = `NOC_X_WIDTH'd2;
    dest_y = `NOC_Y_WIDTH'd20;
end

32'd643:
begin
    dest_x = `NOC_X_WIDTH'd3;
    dest_y = `NOC_Y_WIDTH'd20;
end

32'd644:
begin
    dest_x = `NOC_X_WIDTH'd4;
    dest_y = `NOC_Y_WIDTH'd20;
end

32'd645:
begin
    dest_x = `NOC_X_WIDTH'd5;
    dest_y = `NOC_Y_WIDTH'd20;
end

32'd646:
begin
    dest_x = `NOC_X_WIDTH'd6;
    dest_y = `NOC_Y_WIDTH'd20;
end

32'd647:
begin
    dest_x = `NOC_X_WIDTH'd7;
    dest_y = `NOC_Y_WIDTH'd20;
end

32'd648:
begin
    dest_x = `NOC_X_WIDTH'd8;
    dest_y = `NOC_Y_WIDTH'd20;
end

32'd649:
begin
    dest_x = `NOC_X_WIDTH'd9;
    dest_y = `NOC_Y_WIDTH'd20;
end

32'd650:
begin
    dest_x = `NOC_X_WIDTH'd10;
    dest_y = `NOC_Y_WIDTH'd20;
end

32'd651:
begin
    dest_x = `NOC_X_WIDTH'd11;
    dest_y = `NOC_Y_WIDTH'd20;
end

32'd652:
begin
    dest_x = `NOC_X_WIDTH'd12;
    dest_y = `NOC_Y_WIDTH'd20;
end

32'd653:
begin
    dest_x = `NOC_X_WIDTH'd13;
    dest_y = `NOC_Y_WIDTH'd20;
end

32'd654:
begin
    dest_x = `NOC_X_WIDTH'd14;
    dest_y = `NOC_Y_WIDTH'd20;
end

32'd655:
begin
    dest_x = `NOC_X_WIDTH'd15;
    dest_y = `NOC_Y_WIDTH'd20;
end

32'd656:
begin
    dest_x = `NOC_X_WIDTH'd16;
    dest_y = `NOC_Y_WIDTH'd20;
end

32'd657:
begin
    dest_x = `NOC_X_WIDTH'd17;
    dest_y = `NOC_Y_WIDTH'd20;
end

32'd658:
begin
    dest_x = `NOC_X_WIDTH'd18;
    dest_y = `NOC_Y_WIDTH'd20;
end

32'd659:
begin
    dest_x = `NOC_X_WIDTH'd19;
    dest_y = `NOC_Y_WIDTH'd20;
end

32'd660:
begin
    dest_x = `NOC_X_WIDTH'd20;
    dest_y = `NOC_Y_WIDTH'd20;
end

32'd661:
begin
    dest_x = `NOC_X_WIDTH'd21;
    dest_y = `NOC_Y_WIDTH'd20;
end

32'd662:
begin
    dest_x = `NOC_X_WIDTH'd22;
    dest_y = `NOC_Y_WIDTH'd20;
end

32'd663:
begin
    dest_x = `NOC_X_WIDTH'd23;
    dest_y = `NOC_Y_WIDTH'd20;
end

32'd664:
begin
    dest_x = `NOC_X_WIDTH'd24;
    dest_y = `NOC_Y_WIDTH'd20;
end

32'd665:
begin
    dest_x = `NOC_X_WIDTH'd25;
    dest_y = `NOC_Y_WIDTH'd20;
end

32'd666:
begin
    dest_x = `NOC_X_WIDTH'd26;
    dest_y = `NOC_Y_WIDTH'd20;
end

32'd667:
begin
    dest_x = `NOC_X_WIDTH'd27;
    dest_y = `NOC_Y_WIDTH'd20;
end

32'd668:
begin
    dest_x = `NOC_X_WIDTH'd28;
    dest_y = `NOC_Y_WIDTH'd20;
end

32'd669:
begin
    dest_x = `NOC_X_WIDTH'd29;
    dest_y = `NOC_Y_WIDTH'd20;
end

32'd670:
begin
    dest_x = `NOC_X_WIDTH'd30;
    dest_y = `NOC_Y_WIDTH'd20;
end

32'd671:
begin
    dest_x = `NOC_X_WIDTH'd31;
    dest_y = `NOC_Y_WIDTH'd20;
end

32'd672:
begin
    dest_x = `NOC_X_WIDTH'd0;
    dest_y = `NOC_Y_WIDTH'd21;
end

32'd673:
begin
    dest_x = `NOC_X_WIDTH'd1;
    dest_y = `NOC_Y_WIDTH'd21;
end

32'd674:
begin
    dest_x = `NOC_X_WIDTH'd2;
    dest_y = `NOC_Y_WIDTH'd21;
end

32'd675:
begin
    dest_x = `NOC_X_WIDTH'd3;
    dest_y = `NOC_Y_WIDTH'd21;
end

32'd676:
begin
    dest_x = `NOC_X_WIDTH'd4;
    dest_y = `NOC_Y_WIDTH'd21;
end

32'd677:
begin
    dest_x = `NOC_X_WIDTH'd5;
    dest_y = `NOC_Y_WIDTH'd21;
end

32'd678:
begin
    dest_x = `NOC_X_WIDTH'd6;
    dest_y = `NOC_Y_WIDTH'd21;
end

32'd679:
begin
    dest_x = `NOC_X_WIDTH'd7;
    dest_y = `NOC_Y_WIDTH'd21;
end

32'd680:
begin
    dest_x = `NOC_X_WIDTH'd8;
    dest_y = `NOC_Y_WIDTH'd21;
end

32'd681:
begin
    dest_x = `NOC_X_WIDTH'd9;
    dest_y = `NOC_Y_WIDTH'd21;
end

32'd682:
begin
    dest_x = `NOC_X_WIDTH'd10;
    dest_y = `NOC_Y_WIDTH'd21;
end

32'd683:
begin
    dest_x = `NOC_X_WIDTH'd11;
    dest_y = `NOC_Y_WIDTH'd21;
end

32'd684:
begin
    dest_x = `NOC_X_WIDTH'd12;
    dest_y = `NOC_Y_WIDTH'd21;
end

32'd685:
begin
    dest_x = `NOC_X_WIDTH'd13;
    dest_y = `NOC_Y_WIDTH'd21;
end

32'd686:
begin
    dest_x = `NOC_X_WIDTH'd14;
    dest_y = `NOC_Y_WIDTH'd21;
end

32'd687:
begin
    dest_x = `NOC_X_WIDTH'd15;
    dest_y = `NOC_Y_WIDTH'd21;
end

32'd688:
begin
    dest_x = `NOC_X_WIDTH'd16;
    dest_y = `NOC_Y_WIDTH'd21;
end

32'd689:
begin
    dest_x = `NOC_X_WIDTH'd17;
    dest_y = `NOC_Y_WIDTH'd21;
end

32'd690:
begin
    dest_x = `NOC_X_WIDTH'd18;
    dest_y = `NOC_Y_WIDTH'd21;
end

32'd691:
begin
    dest_x = `NOC_X_WIDTH'd19;
    dest_y = `NOC_Y_WIDTH'd21;
end

32'd692:
begin
    dest_x = `NOC_X_WIDTH'd20;
    dest_y = `NOC_Y_WIDTH'd21;
end

32'd693:
begin
    dest_x = `NOC_X_WIDTH'd21;
    dest_y = `NOC_Y_WIDTH'd21;
end

32'd694:
begin
    dest_x = `NOC_X_WIDTH'd22;
    dest_y = `NOC_Y_WIDTH'd21;
end

32'd695:
begin
    dest_x = `NOC_X_WIDTH'd23;
    dest_y = `NOC_Y_WIDTH'd21;
end

32'd696:
begin
    dest_x = `NOC_X_WIDTH'd24;
    dest_y = `NOC_Y_WIDTH'd21;
end

32'd697:
begin
    dest_x = `NOC_X_WIDTH'd25;
    dest_y = `NOC_Y_WIDTH'd21;
end

32'd698:
begin
    dest_x = `NOC_X_WIDTH'd26;
    dest_y = `NOC_Y_WIDTH'd21;
end

32'd699:
begin
    dest_x = `NOC_X_WIDTH'd27;
    dest_y = `NOC_Y_WIDTH'd21;
end

32'd700:
begin
    dest_x = `NOC_X_WIDTH'd28;
    dest_y = `NOC_Y_WIDTH'd21;
end

32'd701:
begin
    dest_x = `NOC_X_WIDTH'd29;
    dest_y = `NOC_Y_WIDTH'd21;
end

32'd702:
begin
    dest_x = `NOC_X_WIDTH'd30;
    dest_y = `NOC_Y_WIDTH'd21;
end

32'd703:
begin
    dest_x = `NOC_X_WIDTH'd31;
    dest_y = `NOC_Y_WIDTH'd21;
end

32'd704:
begin
    dest_x = `NOC_X_WIDTH'd0;
    dest_y = `NOC_Y_WIDTH'd22;
end

32'd705:
begin
    dest_x = `NOC_X_WIDTH'd1;
    dest_y = `NOC_Y_WIDTH'd22;
end

32'd706:
begin
    dest_x = `NOC_X_WIDTH'd2;
    dest_y = `NOC_Y_WIDTH'd22;
end

32'd707:
begin
    dest_x = `NOC_X_WIDTH'd3;
    dest_y = `NOC_Y_WIDTH'd22;
end

32'd708:
begin
    dest_x = `NOC_X_WIDTH'd4;
    dest_y = `NOC_Y_WIDTH'd22;
end

32'd709:
begin
    dest_x = `NOC_X_WIDTH'd5;
    dest_y = `NOC_Y_WIDTH'd22;
end

32'd710:
begin
    dest_x = `NOC_X_WIDTH'd6;
    dest_y = `NOC_Y_WIDTH'd22;
end

32'd711:
begin
    dest_x = `NOC_X_WIDTH'd7;
    dest_y = `NOC_Y_WIDTH'd22;
end

32'd712:
begin
    dest_x = `NOC_X_WIDTH'd8;
    dest_y = `NOC_Y_WIDTH'd22;
end

32'd713:
begin
    dest_x = `NOC_X_WIDTH'd9;
    dest_y = `NOC_Y_WIDTH'd22;
end

32'd714:
begin
    dest_x = `NOC_X_WIDTH'd10;
    dest_y = `NOC_Y_WIDTH'd22;
end

32'd715:
begin
    dest_x = `NOC_X_WIDTH'd11;
    dest_y = `NOC_Y_WIDTH'd22;
end

32'd716:
begin
    dest_x = `NOC_X_WIDTH'd12;
    dest_y = `NOC_Y_WIDTH'd22;
end

32'd717:
begin
    dest_x = `NOC_X_WIDTH'd13;
    dest_y = `NOC_Y_WIDTH'd22;
end

32'd718:
begin
    dest_x = `NOC_X_WIDTH'd14;
    dest_y = `NOC_Y_WIDTH'd22;
end

32'd719:
begin
    dest_x = `NOC_X_WIDTH'd15;
    dest_y = `NOC_Y_WIDTH'd22;
end

32'd720:
begin
    dest_x = `NOC_X_WIDTH'd16;
    dest_y = `NOC_Y_WIDTH'd22;
end

32'd721:
begin
    dest_x = `NOC_X_WIDTH'd17;
    dest_y = `NOC_Y_WIDTH'd22;
end

32'd722:
begin
    dest_x = `NOC_X_WIDTH'd18;
    dest_y = `NOC_Y_WIDTH'd22;
end

32'd723:
begin
    dest_x = `NOC_X_WIDTH'd19;
    dest_y = `NOC_Y_WIDTH'd22;
end

32'd724:
begin
    dest_x = `NOC_X_WIDTH'd20;
    dest_y = `NOC_Y_WIDTH'd22;
end

32'd725:
begin
    dest_x = `NOC_X_WIDTH'd21;
    dest_y = `NOC_Y_WIDTH'd22;
end

32'd726:
begin
    dest_x = `NOC_X_WIDTH'd22;
    dest_y = `NOC_Y_WIDTH'd22;
end

32'd727:
begin
    dest_x = `NOC_X_WIDTH'd23;
    dest_y = `NOC_Y_WIDTH'd22;
end

32'd728:
begin
    dest_x = `NOC_X_WIDTH'd24;
    dest_y = `NOC_Y_WIDTH'd22;
end

32'd729:
begin
    dest_x = `NOC_X_WIDTH'd25;
    dest_y = `NOC_Y_WIDTH'd22;
end

32'd730:
begin
    dest_x = `NOC_X_WIDTH'd26;
    dest_y = `NOC_Y_WIDTH'd22;
end

32'd731:
begin
    dest_x = `NOC_X_WIDTH'd27;
    dest_y = `NOC_Y_WIDTH'd22;
end

32'd732:
begin
    dest_x = `NOC_X_WIDTH'd28;
    dest_y = `NOC_Y_WIDTH'd22;
end

32'd733:
begin
    dest_x = `NOC_X_WIDTH'd29;
    dest_y = `NOC_Y_WIDTH'd22;
end

32'd734:
begin
    dest_x = `NOC_X_WIDTH'd30;
    dest_y = `NOC_Y_WIDTH'd22;
end

32'd735:
begin
    dest_x = `NOC_X_WIDTH'd31;
    dest_y = `NOC_Y_WIDTH'd22;
end

32'd736:
begin
    dest_x = `NOC_X_WIDTH'd0;
    dest_y = `NOC_Y_WIDTH'd23;
end

32'd737:
begin
    dest_x = `NOC_X_WIDTH'd1;
    dest_y = `NOC_Y_WIDTH'd23;
end

32'd738:
begin
    dest_x = `NOC_X_WIDTH'd2;
    dest_y = `NOC_Y_WIDTH'd23;
end

32'd739:
begin
    dest_x = `NOC_X_WIDTH'd3;
    dest_y = `NOC_Y_WIDTH'd23;
end

32'd740:
begin
    dest_x = `NOC_X_WIDTH'd4;
    dest_y = `NOC_Y_WIDTH'd23;
end

32'd741:
begin
    dest_x = `NOC_X_WIDTH'd5;
    dest_y = `NOC_Y_WIDTH'd23;
end

32'd742:
begin
    dest_x = `NOC_X_WIDTH'd6;
    dest_y = `NOC_Y_WIDTH'd23;
end

32'd743:
begin
    dest_x = `NOC_X_WIDTH'd7;
    dest_y = `NOC_Y_WIDTH'd23;
end

32'd744:
begin
    dest_x = `NOC_X_WIDTH'd8;
    dest_y = `NOC_Y_WIDTH'd23;
end

32'd745:
begin
    dest_x = `NOC_X_WIDTH'd9;
    dest_y = `NOC_Y_WIDTH'd23;
end

32'd746:
begin
    dest_x = `NOC_X_WIDTH'd10;
    dest_y = `NOC_Y_WIDTH'd23;
end

32'd747:
begin
    dest_x = `NOC_X_WIDTH'd11;
    dest_y = `NOC_Y_WIDTH'd23;
end

32'd748:
begin
    dest_x = `NOC_X_WIDTH'd12;
    dest_y = `NOC_Y_WIDTH'd23;
end

32'd749:
begin
    dest_x = `NOC_X_WIDTH'd13;
    dest_y = `NOC_Y_WIDTH'd23;
end

32'd750:
begin
    dest_x = `NOC_X_WIDTH'd14;
    dest_y = `NOC_Y_WIDTH'd23;
end

32'd751:
begin
    dest_x = `NOC_X_WIDTH'd15;
    dest_y = `NOC_Y_WIDTH'd23;
end

32'd752:
begin
    dest_x = `NOC_X_WIDTH'd16;
    dest_y = `NOC_Y_WIDTH'd23;
end

32'd753:
begin
    dest_x = `NOC_X_WIDTH'd17;
    dest_y = `NOC_Y_WIDTH'd23;
end

32'd754:
begin
    dest_x = `NOC_X_WIDTH'd18;
    dest_y = `NOC_Y_WIDTH'd23;
end

32'd755:
begin
    dest_x = `NOC_X_WIDTH'd19;
    dest_y = `NOC_Y_WIDTH'd23;
end

32'd756:
begin
    dest_x = `NOC_X_WIDTH'd20;
    dest_y = `NOC_Y_WIDTH'd23;
end

32'd757:
begin
    dest_x = `NOC_X_WIDTH'd21;
    dest_y = `NOC_Y_WIDTH'd23;
end

32'd758:
begin
    dest_x = `NOC_X_WIDTH'd22;
    dest_y = `NOC_Y_WIDTH'd23;
end

32'd759:
begin
    dest_x = `NOC_X_WIDTH'd23;
    dest_y = `NOC_Y_WIDTH'd23;
end

32'd760:
begin
    dest_x = `NOC_X_WIDTH'd24;
    dest_y = `NOC_Y_WIDTH'd23;
end

32'd761:
begin
    dest_x = `NOC_X_WIDTH'd25;
    dest_y = `NOC_Y_WIDTH'd23;
end

32'd762:
begin
    dest_x = `NOC_X_WIDTH'd26;
    dest_y = `NOC_Y_WIDTH'd23;
end

32'd763:
begin
    dest_x = `NOC_X_WIDTH'd27;
    dest_y = `NOC_Y_WIDTH'd23;
end

32'd764:
begin
    dest_x = `NOC_X_WIDTH'd28;
    dest_y = `NOC_Y_WIDTH'd23;
end

32'd765:
begin
    dest_x = `NOC_X_WIDTH'd29;
    dest_y = `NOC_Y_WIDTH'd23;
end

32'd766:
begin
    dest_x = `NOC_X_WIDTH'd30;
    dest_y = `NOC_Y_WIDTH'd23;
end

32'd767:
begin
    dest_x = `NOC_X_WIDTH'd31;
    dest_y = `NOC_Y_WIDTH'd23;
end

32'd768:
begin
    dest_x = `NOC_X_WIDTH'd0;
    dest_y = `NOC_Y_WIDTH'd24;
end

32'd769:
begin
    dest_x = `NOC_X_WIDTH'd1;
    dest_y = `NOC_Y_WIDTH'd24;
end

32'd770:
begin
    dest_x = `NOC_X_WIDTH'd2;
    dest_y = `NOC_Y_WIDTH'd24;
end

32'd771:
begin
    dest_x = `NOC_X_WIDTH'd3;
    dest_y = `NOC_Y_WIDTH'd24;
end

32'd772:
begin
    dest_x = `NOC_X_WIDTH'd4;
    dest_y = `NOC_Y_WIDTH'd24;
end

32'd773:
begin
    dest_x = `NOC_X_WIDTH'd5;
    dest_y = `NOC_Y_WIDTH'd24;
end

32'd774:
begin
    dest_x = `NOC_X_WIDTH'd6;
    dest_y = `NOC_Y_WIDTH'd24;
end

32'd775:
begin
    dest_x = `NOC_X_WIDTH'd7;
    dest_y = `NOC_Y_WIDTH'd24;
end

32'd776:
begin
    dest_x = `NOC_X_WIDTH'd8;
    dest_y = `NOC_Y_WIDTH'd24;
end

32'd777:
begin
    dest_x = `NOC_X_WIDTH'd9;
    dest_y = `NOC_Y_WIDTH'd24;
end

32'd778:
begin
    dest_x = `NOC_X_WIDTH'd10;
    dest_y = `NOC_Y_WIDTH'd24;
end

32'd779:
begin
    dest_x = `NOC_X_WIDTH'd11;
    dest_y = `NOC_Y_WIDTH'd24;
end

32'd780:
begin
    dest_x = `NOC_X_WIDTH'd12;
    dest_y = `NOC_Y_WIDTH'd24;
end

32'd781:
begin
    dest_x = `NOC_X_WIDTH'd13;
    dest_y = `NOC_Y_WIDTH'd24;
end

32'd782:
begin
    dest_x = `NOC_X_WIDTH'd14;
    dest_y = `NOC_Y_WIDTH'd24;
end

32'd783:
begin
    dest_x = `NOC_X_WIDTH'd15;
    dest_y = `NOC_Y_WIDTH'd24;
end

32'd784:
begin
    dest_x = `NOC_X_WIDTH'd16;
    dest_y = `NOC_Y_WIDTH'd24;
end

32'd785:
begin
    dest_x = `NOC_X_WIDTH'd17;
    dest_y = `NOC_Y_WIDTH'd24;
end

32'd786:
begin
    dest_x = `NOC_X_WIDTH'd18;
    dest_y = `NOC_Y_WIDTH'd24;
end

32'd787:
begin
    dest_x = `NOC_X_WIDTH'd19;
    dest_y = `NOC_Y_WIDTH'd24;
end

32'd788:
begin
    dest_x = `NOC_X_WIDTH'd20;
    dest_y = `NOC_Y_WIDTH'd24;
end

32'd789:
begin
    dest_x = `NOC_X_WIDTH'd21;
    dest_y = `NOC_Y_WIDTH'd24;
end

32'd790:
begin
    dest_x = `NOC_X_WIDTH'd22;
    dest_y = `NOC_Y_WIDTH'd24;
end

32'd791:
begin
    dest_x = `NOC_X_WIDTH'd23;
    dest_y = `NOC_Y_WIDTH'd24;
end

32'd792:
begin
    dest_x = `NOC_X_WIDTH'd24;
    dest_y = `NOC_Y_WIDTH'd24;
end

32'd793:
begin
    dest_x = `NOC_X_WIDTH'd25;
    dest_y = `NOC_Y_WIDTH'd24;
end

32'd794:
begin
    dest_x = `NOC_X_WIDTH'd26;
    dest_y = `NOC_Y_WIDTH'd24;
end

32'd795:
begin
    dest_x = `NOC_X_WIDTH'd27;
    dest_y = `NOC_Y_WIDTH'd24;
end

32'd796:
begin
    dest_x = `NOC_X_WIDTH'd28;
    dest_y = `NOC_Y_WIDTH'd24;
end

32'd797:
begin
    dest_x = `NOC_X_WIDTH'd29;
    dest_y = `NOC_Y_WIDTH'd24;
end

32'd798:
begin
    dest_x = `NOC_X_WIDTH'd30;
    dest_y = `NOC_Y_WIDTH'd24;
end

32'd799:
begin
    dest_x = `NOC_X_WIDTH'd31;
    dest_y = `NOC_Y_WIDTH'd24;
end

32'd800:
begin
    dest_x = `NOC_X_WIDTH'd0;
    dest_y = `NOC_Y_WIDTH'd25;
end

32'd801:
begin
    dest_x = `NOC_X_WIDTH'd1;
    dest_y = `NOC_Y_WIDTH'd25;
end

32'd802:
begin
    dest_x = `NOC_X_WIDTH'd2;
    dest_y = `NOC_Y_WIDTH'd25;
end

32'd803:
begin
    dest_x = `NOC_X_WIDTH'd3;
    dest_y = `NOC_Y_WIDTH'd25;
end

32'd804:
begin
    dest_x = `NOC_X_WIDTH'd4;
    dest_y = `NOC_Y_WIDTH'd25;
end

32'd805:
begin
    dest_x = `NOC_X_WIDTH'd5;
    dest_y = `NOC_Y_WIDTH'd25;
end

32'd806:
begin
    dest_x = `NOC_X_WIDTH'd6;
    dest_y = `NOC_Y_WIDTH'd25;
end

32'd807:
begin
    dest_x = `NOC_X_WIDTH'd7;
    dest_y = `NOC_Y_WIDTH'd25;
end

32'd808:
begin
    dest_x = `NOC_X_WIDTH'd8;
    dest_y = `NOC_Y_WIDTH'd25;
end

32'd809:
begin
    dest_x = `NOC_X_WIDTH'd9;
    dest_y = `NOC_Y_WIDTH'd25;
end

32'd810:
begin
    dest_x = `NOC_X_WIDTH'd10;
    dest_y = `NOC_Y_WIDTH'd25;
end

32'd811:
begin
    dest_x = `NOC_X_WIDTH'd11;
    dest_y = `NOC_Y_WIDTH'd25;
end

32'd812:
begin
    dest_x = `NOC_X_WIDTH'd12;
    dest_y = `NOC_Y_WIDTH'd25;
end

32'd813:
begin
    dest_x = `NOC_X_WIDTH'd13;
    dest_y = `NOC_Y_WIDTH'd25;
end

32'd814:
begin
    dest_x = `NOC_X_WIDTH'd14;
    dest_y = `NOC_Y_WIDTH'd25;
end

32'd815:
begin
    dest_x = `NOC_X_WIDTH'd15;
    dest_y = `NOC_Y_WIDTH'd25;
end

32'd816:
begin
    dest_x = `NOC_X_WIDTH'd16;
    dest_y = `NOC_Y_WIDTH'd25;
end

32'd817:
begin
    dest_x = `NOC_X_WIDTH'd17;
    dest_y = `NOC_Y_WIDTH'd25;
end

32'd818:
begin
    dest_x = `NOC_X_WIDTH'd18;
    dest_y = `NOC_Y_WIDTH'd25;
end

32'd819:
begin
    dest_x = `NOC_X_WIDTH'd19;
    dest_y = `NOC_Y_WIDTH'd25;
end

32'd820:
begin
    dest_x = `NOC_X_WIDTH'd20;
    dest_y = `NOC_Y_WIDTH'd25;
end

32'd821:
begin
    dest_x = `NOC_X_WIDTH'd21;
    dest_y = `NOC_Y_WIDTH'd25;
end

32'd822:
begin
    dest_x = `NOC_X_WIDTH'd22;
    dest_y = `NOC_Y_WIDTH'd25;
end

32'd823:
begin
    dest_x = `NOC_X_WIDTH'd23;
    dest_y = `NOC_Y_WIDTH'd25;
end

32'd824:
begin
    dest_x = `NOC_X_WIDTH'd24;
    dest_y = `NOC_Y_WIDTH'd25;
end

32'd825:
begin
    dest_x = `NOC_X_WIDTH'd25;
    dest_y = `NOC_Y_WIDTH'd25;
end

32'd826:
begin
    dest_x = `NOC_X_WIDTH'd26;
    dest_y = `NOC_Y_WIDTH'd25;
end

32'd827:
begin
    dest_x = `NOC_X_WIDTH'd27;
    dest_y = `NOC_Y_WIDTH'd25;
end

32'd828:
begin
    dest_x = `NOC_X_WIDTH'd28;
    dest_y = `NOC_Y_WIDTH'd25;
end

32'd829:
begin
    dest_x = `NOC_X_WIDTH'd29;
    dest_y = `NOC_Y_WIDTH'd25;
end

32'd830:
begin
    dest_x = `NOC_X_WIDTH'd30;
    dest_y = `NOC_Y_WIDTH'd25;
end

32'd831:
begin
    dest_x = `NOC_X_WIDTH'd31;
    dest_y = `NOC_Y_WIDTH'd25;
end

32'd832:
begin
    dest_x = `NOC_X_WIDTH'd0;
    dest_y = `NOC_Y_WIDTH'd26;
end

32'd833:
begin
    dest_x = `NOC_X_WIDTH'd1;
    dest_y = `NOC_Y_WIDTH'd26;
end

32'd834:
begin
    dest_x = `NOC_X_WIDTH'd2;
    dest_y = `NOC_Y_WIDTH'd26;
end

32'd835:
begin
    dest_x = `NOC_X_WIDTH'd3;
    dest_y = `NOC_Y_WIDTH'd26;
end

32'd836:
begin
    dest_x = `NOC_X_WIDTH'd4;
    dest_y = `NOC_Y_WIDTH'd26;
end

32'd837:
begin
    dest_x = `NOC_X_WIDTH'd5;
    dest_y = `NOC_Y_WIDTH'd26;
end

32'd838:
begin
    dest_x = `NOC_X_WIDTH'd6;
    dest_y = `NOC_Y_WIDTH'd26;
end

32'd839:
begin
    dest_x = `NOC_X_WIDTH'd7;
    dest_y = `NOC_Y_WIDTH'd26;
end

32'd840:
begin
    dest_x = `NOC_X_WIDTH'd8;
    dest_y = `NOC_Y_WIDTH'd26;
end

32'd841:
begin
    dest_x = `NOC_X_WIDTH'd9;
    dest_y = `NOC_Y_WIDTH'd26;
end

32'd842:
begin
    dest_x = `NOC_X_WIDTH'd10;
    dest_y = `NOC_Y_WIDTH'd26;
end

32'd843:
begin
    dest_x = `NOC_X_WIDTH'd11;
    dest_y = `NOC_Y_WIDTH'd26;
end

32'd844:
begin
    dest_x = `NOC_X_WIDTH'd12;
    dest_y = `NOC_Y_WIDTH'd26;
end

32'd845:
begin
    dest_x = `NOC_X_WIDTH'd13;
    dest_y = `NOC_Y_WIDTH'd26;
end

32'd846:
begin
    dest_x = `NOC_X_WIDTH'd14;
    dest_y = `NOC_Y_WIDTH'd26;
end

32'd847:
begin
    dest_x = `NOC_X_WIDTH'd15;
    dest_y = `NOC_Y_WIDTH'd26;
end

32'd848:
begin
    dest_x = `NOC_X_WIDTH'd16;
    dest_y = `NOC_Y_WIDTH'd26;
end

32'd849:
begin
    dest_x = `NOC_X_WIDTH'd17;
    dest_y = `NOC_Y_WIDTH'd26;
end

32'd850:
begin
    dest_x = `NOC_X_WIDTH'd18;
    dest_y = `NOC_Y_WIDTH'd26;
end

32'd851:
begin
    dest_x = `NOC_X_WIDTH'd19;
    dest_y = `NOC_Y_WIDTH'd26;
end

32'd852:
begin
    dest_x = `NOC_X_WIDTH'd20;
    dest_y = `NOC_Y_WIDTH'd26;
end

32'd853:
begin
    dest_x = `NOC_X_WIDTH'd21;
    dest_y = `NOC_Y_WIDTH'd26;
end

32'd854:
begin
    dest_x = `NOC_X_WIDTH'd22;
    dest_y = `NOC_Y_WIDTH'd26;
end

32'd855:
begin
    dest_x = `NOC_X_WIDTH'd23;
    dest_y = `NOC_Y_WIDTH'd26;
end

32'd856:
begin
    dest_x = `NOC_X_WIDTH'd24;
    dest_y = `NOC_Y_WIDTH'd26;
end

32'd857:
begin
    dest_x = `NOC_X_WIDTH'd25;
    dest_y = `NOC_Y_WIDTH'd26;
end

32'd858:
begin
    dest_x = `NOC_X_WIDTH'd26;
    dest_y = `NOC_Y_WIDTH'd26;
end

32'd859:
begin
    dest_x = `NOC_X_WIDTH'd27;
    dest_y = `NOC_Y_WIDTH'd26;
end

32'd860:
begin
    dest_x = `NOC_X_WIDTH'd28;
    dest_y = `NOC_Y_WIDTH'd26;
end

32'd861:
begin
    dest_x = `NOC_X_WIDTH'd29;
    dest_y = `NOC_Y_WIDTH'd26;
end

32'd862:
begin
    dest_x = `NOC_X_WIDTH'd30;
    dest_y = `NOC_Y_WIDTH'd26;
end

32'd863:
begin
    dest_x = `NOC_X_WIDTH'd31;
    dest_y = `NOC_Y_WIDTH'd26;
end

32'd864:
begin
    dest_x = `NOC_X_WIDTH'd0;
    dest_y = `NOC_Y_WIDTH'd27;
end

32'd865:
begin
    dest_x = `NOC_X_WIDTH'd1;
    dest_y = `NOC_Y_WIDTH'd27;
end

32'd866:
begin
    dest_x = `NOC_X_WIDTH'd2;
    dest_y = `NOC_Y_WIDTH'd27;
end

32'd867:
begin
    dest_x = `NOC_X_WIDTH'd3;
    dest_y = `NOC_Y_WIDTH'd27;
end

32'd868:
begin
    dest_x = `NOC_X_WIDTH'd4;
    dest_y = `NOC_Y_WIDTH'd27;
end

32'd869:
begin
    dest_x = `NOC_X_WIDTH'd5;
    dest_y = `NOC_Y_WIDTH'd27;
end

32'd870:
begin
    dest_x = `NOC_X_WIDTH'd6;
    dest_y = `NOC_Y_WIDTH'd27;
end

32'd871:
begin
    dest_x = `NOC_X_WIDTH'd7;
    dest_y = `NOC_Y_WIDTH'd27;
end

32'd872:
begin
    dest_x = `NOC_X_WIDTH'd8;
    dest_y = `NOC_Y_WIDTH'd27;
end

32'd873:
begin
    dest_x = `NOC_X_WIDTH'd9;
    dest_y = `NOC_Y_WIDTH'd27;
end

32'd874:
begin
    dest_x = `NOC_X_WIDTH'd10;
    dest_y = `NOC_Y_WIDTH'd27;
end

32'd875:
begin
    dest_x = `NOC_X_WIDTH'd11;
    dest_y = `NOC_Y_WIDTH'd27;
end

32'd876:
begin
    dest_x = `NOC_X_WIDTH'd12;
    dest_y = `NOC_Y_WIDTH'd27;
end

32'd877:
begin
    dest_x = `NOC_X_WIDTH'd13;
    dest_y = `NOC_Y_WIDTH'd27;
end

32'd878:
begin
    dest_x = `NOC_X_WIDTH'd14;
    dest_y = `NOC_Y_WIDTH'd27;
end

32'd879:
begin
    dest_x = `NOC_X_WIDTH'd15;
    dest_y = `NOC_Y_WIDTH'd27;
end

32'd880:
begin
    dest_x = `NOC_X_WIDTH'd16;
    dest_y = `NOC_Y_WIDTH'd27;
end

32'd881:
begin
    dest_x = `NOC_X_WIDTH'd17;
    dest_y = `NOC_Y_WIDTH'd27;
end

32'd882:
begin
    dest_x = `NOC_X_WIDTH'd18;
    dest_y = `NOC_Y_WIDTH'd27;
end

32'd883:
begin
    dest_x = `NOC_X_WIDTH'd19;
    dest_y = `NOC_Y_WIDTH'd27;
end

32'd884:
begin
    dest_x = `NOC_X_WIDTH'd20;
    dest_y = `NOC_Y_WIDTH'd27;
end

32'd885:
begin
    dest_x = `NOC_X_WIDTH'd21;
    dest_y = `NOC_Y_WIDTH'd27;
end

32'd886:
begin
    dest_x = `NOC_X_WIDTH'd22;
    dest_y = `NOC_Y_WIDTH'd27;
end

32'd887:
begin
    dest_x = `NOC_X_WIDTH'd23;
    dest_y = `NOC_Y_WIDTH'd27;
end

32'd888:
begin
    dest_x = `NOC_X_WIDTH'd24;
    dest_y = `NOC_Y_WIDTH'd27;
end

32'd889:
begin
    dest_x = `NOC_X_WIDTH'd25;
    dest_y = `NOC_Y_WIDTH'd27;
end

32'd890:
begin
    dest_x = `NOC_X_WIDTH'd26;
    dest_y = `NOC_Y_WIDTH'd27;
end

32'd891:
begin
    dest_x = `NOC_X_WIDTH'd27;
    dest_y = `NOC_Y_WIDTH'd27;
end

32'd892:
begin
    dest_x = `NOC_X_WIDTH'd28;
    dest_y = `NOC_Y_WIDTH'd27;
end

32'd893:
begin
    dest_x = `NOC_X_WIDTH'd29;
    dest_y = `NOC_Y_WIDTH'd27;
end

32'd894:
begin
    dest_x = `NOC_X_WIDTH'd30;
    dest_y = `NOC_Y_WIDTH'd27;
end

32'd895:
begin
    dest_x = `NOC_X_WIDTH'd31;
    dest_y = `NOC_Y_WIDTH'd27;
end

32'd896:
begin
    dest_x = `NOC_X_WIDTH'd0;
    dest_y = `NOC_Y_WIDTH'd28;
end

32'd897:
begin
    dest_x = `NOC_X_WIDTH'd1;
    dest_y = `NOC_Y_WIDTH'd28;
end

32'd898:
begin
    dest_x = `NOC_X_WIDTH'd2;
    dest_y = `NOC_Y_WIDTH'd28;
end

32'd899:
begin
    dest_x = `NOC_X_WIDTH'd3;
    dest_y = `NOC_Y_WIDTH'd28;
end

32'd900:
begin
    dest_x = `NOC_X_WIDTH'd4;
    dest_y = `NOC_Y_WIDTH'd28;
end

32'd901:
begin
    dest_x = `NOC_X_WIDTH'd5;
    dest_y = `NOC_Y_WIDTH'd28;
end

32'd902:
begin
    dest_x = `NOC_X_WIDTH'd6;
    dest_y = `NOC_Y_WIDTH'd28;
end

32'd903:
begin
    dest_x = `NOC_X_WIDTH'd7;
    dest_y = `NOC_Y_WIDTH'd28;
end

32'd904:
begin
    dest_x = `NOC_X_WIDTH'd8;
    dest_y = `NOC_Y_WIDTH'd28;
end

32'd905:
begin
    dest_x = `NOC_X_WIDTH'd9;
    dest_y = `NOC_Y_WIDTH'd28;
end

32'd906:
begin
    dest_x = `NOC_X_WIDTH'd10;
    dest_y = `NOC_Y_WIDTH'd28;
end

32'd907:
begin
    dest_x = `NOC_X_WIDTH'd11;
    dest_y = `NOC_Y_WIDTH'd28;
end

32'd908:
begin
    dest_x = `NOC_X_WIDTH'd12;
    dest_y = `NOC_Y_WIDTH'd28;
end

32'd909:
begin
    dest_x = `NOC_X_WIDTH'd13;
    dest_y = `NOC_Y_WIDTH'd28;
end

32'd910:
begin
    dest_x = `NOC_X_WIDTH'd14;
    dest_y = `NOC_Y_WIDTH'd28;
end

32'd911:
begin
    dest_x = `NOC_X_WIDTH'd15;
    dest_y = `NOC_Y_WIDTH'd28;
end

32'd912:
begin
    dest_x = `NOC_X_WIDTH'd16;
    dest_y = `NOC_Y_WIDTH'd28;
end

32'd913:
begin
    dest_x = `NOC_X_WIDTH'd17;
    dest_y = `NOC_Y_WIDTH'd28;
end

32'd914:
begin
    dest_x = `NOC_X_WIDTH'd18;
    dest_y = `NOC_Y_WIDTH'd28;
end

32'd915:
begin
    dest_x = `NOC_X_WIDTH'd19;
    dest_y = `NOC_Y_WIDTH'd28;
end

32'd916:
begin
    dest_x = `NOC_X_WIDTH'd20;
    dest_y = `NOC_Y_WIDTH'd28;
end

32'd917:
begin
    dest_x = `NOC_X_WIDTH'd21;
    dest_y = `NOC_Y_WIDTH'd28;
end

32'd918:
begin
    dest_x = `NOC_X_WIDTH'd22;
    dest_y = `NOC_Y_WIDTH'd28;
end

32'd919:
begin
    dest_x = `NOC_X_WIDTH'd23;
    dest_y = `NOC_Y_WIDTH'd28;
end

32'd920:
begin
    dest_x = `NOC_X_WIDTH'd24;
    dest_y = `NOC_Y_WIDTH'd28;
end

32'd921:
begin
    dest_x = `NOC_X_WIDTH'd25;
    dest_y = `NOC_Y_WIDTH'd28;
end

32'd922:
begin
    dest_x = `NOC_X_WIDTH'd26;
    dest_y = `NOC_Y_WIDTH'd28;
end

32'd923:
begin
    dest_x = `NOC_X_WIDTH'd27;
    dest_y = `NOC_Y_WIDTH'd28;
end

32'd924:
begin
    dest_x = `NOC_X_WIDTH'd28;
    dest_y = `NOC_Y_WIDTH'd28;
end

32'd925:
begin
    dest_x = `NOC_X_WIDTH'd29;
    dest_y = `NOC_Y_WIDTH'd28;
end

32'd926:
begin
    dest_x = `NOC_X_WIDTH'd30;
    dest_y = `NOC_Y_WIDTH'd28;
end

32'd927:
begin
    dest_x = `NOC_X_WIDTH'd31;
    dest_y = `NOC_Y_WIDTH'd28;
end

32'd928:
begin
    dest_x = `NOC_X_WIDTH'd0;
    dest_y = `NOC_Y_WIDTH'd29;
end

32'd929:
begin
    dest_x = `NOC_X_WIDTH'd1;
    dest_y = `NOC_Y_WIDTH'd29;
end

32'd930:
begin
    dest_x = `NOC_X_WIDTH'd2;
    dest_y = `NOC_Y_WIDTH'd29;
end

32'd931:
begin
    dest_x = `NOC_X_WIDTH'd3;
    dest_y = `NOC_Y_WIDTH'd29;
end

32'd932:
begin
    dest_x = `NOC_X_WIDTH'd4;
    dest_y = `NOC_Y_WIDTH'd29;
end

32'd933:
begin
    dest_x = `NOC_X_WIDTH'd5;
    dest_y = `NOC_Y_WIDTH'd29;
end

32'd934:
begin
    dest_x = `NOC_X_WIDTH'd6;
    dest_y = `NOC_Y_WIDTH'd29;
end

32'd935:
begin
    dest_x = `NOC_X_WIDTH'd7;
    dest_y = `NOC_Y_WIDTH'd29;
end

32'd936:
begin
    dest_x = `NOC_X_WIDTH'd8;
    dest_y = `NOC_Y_WIDTH'd29;
end

32'd937:
begin
    dest_x = `NOC_X_WIDTH'd9;
    dest_y = `NOC_Y_WIDTH'd29;
end

32'd938:
begin
    dest_x = `NOC_X_WIDTH'd10;
    dest_y = `NOC_Y_WIDTH'd29;
end

32'd939:
begin
    dest_x = `NOC_X_WIDTH'd11;
    dest_y = `NOC_Y_WIDTH'd29;
end

32'd940:
begin
    dest_x = `NOC_X_WIDTH'd12;
    dest_y = `NOC_Y_WIDTH'd29;
end

32'd941:
begin
    dest_x = `NOC_X_WIDTH'd13;
    dest_y = `NOC_Y_WIDTH'd29;
end

32'd942:
begin
    dest_x = `NOC_X_WIDTH'd14;
    dest_y = `NOC_Y_WIDTH'd29;
end

32'd943:
begin
    dest_x = `NOC_X_WIDTH'd15;
    dest_y = `NOC_Y_WIDTH'd29;
end

32'd944:
begin
    dest_x = `NOC_X_WIDTH'd16;
    dest_y = `NOC_Y_WIDTH'd29;
end

32'd945:
begin
    dest_x = `NOC_X_WIDTH'd17;
    dest_y = `NOC_Y_WIDTH'd29;
end

32'd946:
begin
    dest_x = `NOC_X_WIDTH'd18;
    dest_y = `NOC_Y_WIDTH'd29;
end

32'd947:
begin
    dest_x = `NOC_X_WIDTH'd19;
    dest_y = `NOC_Y_WIDTH'd29;
end

32'd948:
begin
    dest_x = `NOC_X_WIDTH'd20;
    dest_y = `NOC_Y_WIDTH'd29;
end

32'd949:
begin
    dest_x = `NOC_X_WIDTH'd21;
    dest_y = `NOC_Y_WIDTH'd29;
end

32'd950:
begin
    dest_x = `NOC_X_WIDTH'd22;
    dest_y = `NOC_Y_WIDTH'd29;
end

32'd951:
begin
    dest_x = `NOC_X_WIDTH'd23;
    dest_y = `NOC_Y_WIDTH'd29;
end

32'd952:
begin
    dest_x = `NOC_X_WIDTH'd24;
    dest_y = `NOC_Y_WIDTH'd29;
end

32'd953:
begin
    dest_x = `NOC_X_WIDTH'd25;
    dest_y = `NOC_Y_WIDTH'd29;
end

32'd954:
begin
    dest_x = `NOC_X_WIDTH'd26;
    dest_y = `NOC_Y_WIDTH'd29;
end

32'd955:
begin
    dest_x = `NOC_X_WIDTH'd27;
    dest_y = `NOC_Y_WIDTH'd29;
end

32'd956:
begin
    dest_x = `NOC_X_WIDTH'd28;
    dest_y = `NOC_Y_WIDTH'd29;
end

32'd957:
begin
    dest_x = `NOC_X_WIDTH'd29;
    dest_y = `NOC_Y_WIDTH'd29;
end

32'd958:
begin
    dest_x = `NOC_X_WIDTH'd30;
    dest_y = `NOC_Y_WIDTH'd29;
end

32'd959:
begin
    dest_x = `NOC_X_WIDTH'd31;
    dest_y = `NOC_Y_WIDTH'd29;
end

32'd960:
begin
    dest_x = `NOC_X_WIDTH'd0;
    dest_y = `NOC_Y_WIDTH'd30;
end

32'd961:
begin
    dest_x = `NOC_X_WIDTH'd1;
    dest_y = `NOC_Y_WIDTH'd30;
end

32'd962:
begin
    dest_x = `NOC_X_WIDTH'd2;
    dest_y = `NOC_Y_WIDTH'd30;
end

32'd963:
begin
    dest_x = `NOC_X_WIDTH'd3;
    dest_y = `NOC_Y_WIDTH'd30;
end

32'd964:
begin
    dest_x = `NOC_X_WIDTH'd4;
    dest_y = `NOC_Y_WIDTH'd30;
end

32'd965:
begin
    dest_x = `NOC_X_WIDTH'd5;
    dest_y = `NOC_Y_WIDTH'd30;
end

32'd966:
begin
    dest_x = `NOC_X_WIDTH'd6;
    dest_y = `NOC_Y_WIDTH'd30;
end

32'd967:
begin
    dest_x = `NOC_X_WIDTH'd7;
    dest_y = `NOC_Y_WIDTH'd30;
end

32'd968:
begin
    dest_x = `NOC_X_WIDTH'd8;
    dest_y = `NOC_Y_WIDTH'd30;
end

32'd969:
begin
    dest_x = `NOC_X_WIDTH'd9;
    dest_y = `NOC_Y_WIDTH'd30;
end

32'd970:
begin
    dest_x = `NOC_X_WIDTH'd10;
    dest_y = `NOC_Y_WIDTH'd30;
end

32'd971:
begin
    dest_x = `NOC_X_WIDTH'd11;
    dest_y = `NOC_Y_WIDTH'd30;
end

32'd972:
begin
    dest_x = `NOC_X_WIDTH'd12;
    dest_y = `NOC_Y_WIDTH'd30;
end

32'd973:
begin
    dest_x = `NOC_X_WIDTH'd13;
    dest_y = `NOC_Y_WIDTH'd30;
end

32'd974:
begin
    dest_x = `NOC_X_WIDTH'd14;
    dest_y = `NOC_Y_WIDTH'd30;
end

32'd975:
begin
    dest_x = `NOC_X_WIDTH'd15;
    dest_y = `NOC_Y_WIDTH'd30;
end

32'd976:
begin
    dest_x = `NOC_X_WIDTH'd16;
    dest_y = `NOC_Y_WIDTH'd30;
end

32'd977:
begin
    dest_x = `NOC_X_WIDTH'd17;
    dest_y = `NOC_Y_WIDTH'd30;
end

32'd978:
begin
    dest_x = `NOC_X_WIDTH'd18;
    dest_y = `NOC_Y_WIDTH'd30;
end

32'd979:
begin
    dest_x = `NOC_X_WIDTH'd19;
    dest_y = `NOC_Y_WIDTH'd30;
end

32'd980:
begin
    dest_x = `NOC_X_WIDTH'd20;
    dest_y = `NOC_Y_WIDTH'd30;
end

32'd981:
begin
    dest_x = `NOC_X_WIDTH'd21;
    dest_y = `NOC_Y_WIDTH'd30;
end

32'd982:
begin
    dest_x = `NOC_X_WIDTH'd22;
    dest_y = `NOC_Y_WIDTH'd30;
end

32'd983:
begin
    dest_x = `NOC_X_WIDTH'd23;
    dest_y = `NOC_Y_WIDTH'd30;
end

32'd984:
begin
    dest_x = `NOC_X_WIDTH'd24;
    dest_y = `NOC_Y_WIDTH'd30;
end

32'd985:
begin
    dest_x = `NOC_X_WIDTH'd25;
    dest_y = `NOC_Y_WIDTH'd30;
end

32'd986:
begin
    dest_x = `NOC_X_WIDTH'd26;
    dest_y = `NOC_Y_WIDTH'd30;
end

32'd987:
begin
    dest_x = `NOC_X_WIDTH'd27;
    dest_y = `NOC_Y_WIDTH'd30;
end

32'd988:
begin
    dest_x = `NOC_X_WIDTH'd28;
    dest_y = `NOC_Y_WIDTH'd30;
end

32'd989:
begin
    dest_x = `NOC_X_WIDTH'd29;
    dest_y = `NOC_Y_WIDTH'd30;
end

32'd990:
begin
    dest_x = `NOC_X_WIDTH'd30;
    dest_y = `NOC_Y_WIDTH'd30;
end

32'd991:
begin
    dest_x = `NOC_X_WIDTH'd31;
    dest_y = `NOC_Y_WIDTH'd30;
end

32'd992:
begin
    dest_x = `NOC_X_WIDTH'd0;
    dest_y = `NOC_Y_WIDTH'd31;
end

32'd993:
begin
    dest_x = `NOC_X_WIDTH'd1;
    dest_y = `NOC_Y_WIDTH'd31;
end

32'd994:
begin
    dest_x = `NOC_X_WIDTH'd2;
    dest_y = `NOC_Y_WIDTH'd31;
end

32'd995:
begin
    dest_x = `NOC_X_WIDTH'd3;
    dest_y = `NOC_Y_WIDTH'd31;
end

32'd996:
begin
    dest_x = `NOC_X_WIDTH'd4;
    dest_y = `NOC_Y_WIDTH'd31;
end

32'd997:
begin
    dest_x = `NOC_X_WIDTH'd5;
    dest_y = `NOC_Y_WIDTH'd31;
end

32'd998:
begin
    dest_x = `NOC_X_WIDTH'd6;
    dest_y = `NOC_Y_WIDTH'd31;
end

32'd999:
begin
    dest_x = `NOC_X_WIDTH'd7;
    dest_y = `NOC_Y_WIDTH'd31;
end

32'd1000:
begin
    dest_x = `NOC_X_WIDTH'd8;
    dest_y = `NOC_Y_WIDTH'd31;
end

32'd1001:
begin
    dest_x = `NOC_X_WIDTH'd9;
    dest_y = `NOC_Y_WIDTH'd31;
end

32'd1002:
begin
    dest_x = `NOC_X_WIDTH'd10;
    dest_y = `NOC_Y_WIDTH'd31;
end

32'd1003:
begin
    dest_x = `NOC_X_WIDTH'd11;
    dest_y = `NOC_Y_WIDTH'd31;
end

32'd1004:
begin
    dest_x = `NOC_X_WIDTH'd12;
    dest_y = `NOC_Y_WIDTH'd31;
end

32'd1005:
begin
    dest_x = `NOC_X_WIDTH'd13;
    dest_y = `NOC_Y_WIDTH'd31;
end

32'd1006:
begin
    dest_x = `NOC_X_WIDTH'd14;
    dest_y = `NOC_Y_WIDTH'd31;
end

32'd1007:
begin
    dest_x = `NOC_X_WIDTH'd15;
    dest_y = `NOC_Y_WIDTH'd31;
end

32'd1008:
begin
    dest_x = `NOC_X_WIDTH'd16;
    dest_y = `NOC_Y_WIDTH'd31;
end

32'd1009:
begin
    dest_x = `NOC_X_WIDTH'd17;
    dest_y = `NOC_Y_WIDTH'd31;
end

32'd1010:
begin
    dest_x = `NOC_X_WIDTH'd18;
    dest_y = `NOC_Y_WIDTH'd31;
end

32'd1011:
begin
    dest_x = `NOC_X_WIDTH'd19;
    dest_y = `NOC_Y_WIDTH'd31;
end

32'd1012:
begin
    dest_x = `NOC_X_WIDTH'd20;
    dest_y = `NOC_Y_WIDTH'd31;
end

32'd1013:
begin
    dest_x = `NOC_X_WIDTH'd21;
    dest_y = `NOC_Y_WIDTH'd31;
end

32'd1014:
begin
    dest_x = `NOC_X_WIDTH'd22;
    dest_y = `NOC_Y_WIDTH'd31;
end

32'd1015:
begin
    dest_x = `NOC_X_WIDTH'd23;
    dest_y = `NOC_Y_WIDTH'd31;
end

32'd1016:
begin
    dest_x = `NOC_X_WIDTH'd24;
    dest_y = `NOC_Y_WIDTH'd31;
end

32'd1017:
begin
    dest_x = `NOC_X_WIDTH'd25;
    dest_y = `NOC_Y_WIDTH'd31;
end

32'd1018:
begin
    dest_x = `NOC_X_WIDTH'd26;
    dest_y = `NOC_Y_WIDTH'd31;
end

32'd1019:
begin
    dest_x = `NOC_X_WIDTH'd27;
    dest_y = `NOC_Y_WIDTH'd31;
end

32'd1020:
begin
    dest_x = `NOC_X_WIDTH'd28;
    dest_y = `NOC_Y_WIDTH'd31;
end

32'd1021:
begin
    dest_x = `NOC_X_WIDTH'd29;
    dest_y = `NOC_Y_WIDTH'd31;
end

32'd1022:
begin
    dest_x = `NOC_X_WIDTH'd30;
    dest_y = `NOC_Y_WIDTH'd31;
end

32'd1023:
begin
    dest_x = `NOC_X_WIDTH'd31;
    dest_y = `NOC_Y_WIDTH'd31;
end

    default:
    begin
        dest_x = `NOC_X_WIDTH'dX;
        dest_y = `NOC_Y_WIDTH'dX;
    end
    endcase
end


// input signals

wire                             spc0_inst_done_buf  = spc0_inst_done;
wire [63:0]                      pc_w0_buf           = pc_w0;


wire                             spc1_inst_done_buf  = spc1_inst_done;
wire [63:0]                      pc_w1_buf           = pc_w1;


wire                             spc2_inst_done_buf  = spc2_inst_done;
wire [63:0]                      pc_w2_buf           = pc_w2;


wire                             spc3_inst_done_buf  = spc3_inst_done;
wire [63:0]                      pc_w3_buf           = pc_w3;


wire                             spc4_inst_done_buf  = spc4_inst_done;
wire [63:0]                      pc_w4_buf           = pc_w4;


wire                             spc5_inst_done_buf  = spc5_inst_done;
wire [63:0]                      pc_w5_buf           = pc_w5;


wire                             spc6_inst_done_buf  = spc6_inst_done;
wire [63:0]                      pc_w6_buf           = pc_w6;


wire                             spc7_inst_done_buf  = spc7_inst_done;
wire [63:0]                      pc_w7_buf           = pc_w7;


wire                             spc8_inst_done_buf  = spc8_inst_done;
wire [63:0]                      pc_w8_buf           = pc_w8;


wire                             spc9_inst_done_buf  = spc9_inst_done;
wire [63:0]                      pc_w9_buf           = pc_w9;


wire                             spc10_inst_done_buf  = spc10_inst_done;
wire [63:0]                      pc_w10_buf           = pc_w10;


wire                             spc11_inst_done_buf  = spc11_inst_done;
wire [63:0]                      pc_w11_buf           = pc_w11;


wire                             spc12_inst_done_buf  = spc12_inst_done;
wire [63:0]                      pc_w12_buf           = pc_w12;


wire                             spc13_inst_done_buf  = spc13_inst_done;
wire [63:0]                      pc_w13_buf           = pc_w13;


wire                             spc14_inst_done_buf  = spc14_inst_done;
wire [63:0]                      pc_w14_buf           = pc_w14;


wire                             spc15_inst_done_buf  = spc15_inst_done;
wire [63:0]                      pc_w15_buf           = pc_w15;


wire                             spc16_inst_done_buf  = spc16_inst_done;
wire [63:0]                      pc_w16_buf           = pc_w16;


wire                             spc17_inst_done_buf  = spc17_inst_done;
wire [63:0]                      pc_w17_buf           = pc_w17;


wire                             spc18_inst_done_buf  = spc18_inst_done;
wire [63:0]                      pc_w18_buf           = pc_w18;


wire                             spc19_inst_done_buf  = spc19_inst_done;
wire [63:0]                      pc_w19_buf           = pc_w19;


wire                             spc20_inst_done_buf  = spc20_inst_done;
wire [63:0]                      pc_w20_buf           = pc_w20;


wire                             spc21_inst_done_buf  = spc21_inst_done;
wire [63:0]                      pc_w21_buf           = pc_w21;


wire                             spc22_inst_done_buf  = spc22_inst_done;
wire [63:0]                      pc_w22_buf           = pc_w22;


wire                             spc23_inst_done_buf  = spc23_inst_done;
wire [63:0]                      pc_w23_buf           = pc_w23;


wire                             spc24_inst_done_buf  = spc24_inst_done;
wire [63:0]                      pc_w24_buf           = pc_w24;


wire                             spc25_inst_done_buf  = spc25_inst_done;
wire [63:0]                      pc_w25_buf           = pc_w25;


wire                             spc26_inst_done_buf  = spc26_inst_done;
wire [63:0]                      pc_w26_buf           = pc_w26;


wire                             spc27_inst_done_buf  = spc27_inst_done;
wire [63:0]                      pc_w27_buf           = pc_w27;


wire                             spc28_inst_done_buf  = spc28_inst_done;
wire [63:0]                      pc_w28_buf           = pc_w28;


wire                             spc29_inst_done_buf  = spc29_inst_done;
wire [63:0]                      pc_w29_buf           = pc_w29;


wire                             spc30_inst_done_buf  = spc30_inst_done;
wire [63:0]                      pc_w30_buf           = pc_w30;


wire                             spc31_inst_done_buf  = spc31_inst_done;
wire [63:0]                      pc_w31_buf           = pc_w31;


wire                             spc32_inst_done_buf  = spc32_inst_done;
wire [63:0]                      pc_w32_buf           = pc_w32;


wire                             spc33_inst_done_buf  = spc33_inst_done;
wire [63:0]                      pc_w33_buf           = pc_w33;


wire                             spc34_inst_done_buf  = spc34_inst_done;
wire [63:0]                      pc_w34_buf           = pc_w34;


wire                             spc35_inst_done_buf  = spc35_inst_done;
wire [63:0]                      pc_w35_buf           = pc_w35;


wire                             spc36_inst_done_buf  = spc36_inst_done;
wire [63:0]                      pc_w36_buf           = pc_w36;


wire                             spc37_inst_done_buf  = spc37_inst_done;
wire [63:0]                      pc_w37_buf           = pc_w37;


wire                             spc38_inst_done_buf  = spc38_inst_done;
wire [63:0]                      pc_w38_buf           = pc_w38;


wire                             spc39_inst_done_buf  = spc39_inst_done;
wire [63:0]                      pc_w39_buf           = pc_w39;


wire                             spc40_inst_done_buf  = spc40_inst_done;
wire [63:0]                      pc_w40_buf           = pc_w40;


wire                             spc41_inst_done_buf  = spc41_inst_done;
wire [63:0]                      pc_w41_buf           = pc_w41;


wire                             spc42_inst_done_buf  = spc42_inst_done;
wire [63:0]                      pc_w42_buf           = pc_w42;


wire                             spc43_inst_done_buf  = spc43_inst_done;
wire [63:0]                      pc_w43_buf           = pc_w43;


wire                             spc44_inst_done_buf  = spc44_inst_done;
wire [63:0]                      pc_w44_buf           = pc_w44;


wire                             spc45_inst_done_buf  = spc45_inst_done;
wire [63:0]                      pc_w45_buf           = pc_w45;


wire                             spc46_inst_done_buf  = spc46_inst_done;
wire [63:0]                      pc_w46_buf           = pc_w46;


wire                             spc47_inst_done_buf  = spc47_inst_done;
wire [63:0]                      pc_w47_buf           = pc_w47;


wire                             spc48_inst_done_buf  = spc48_inst_done;
wire [63:0]                      pc_w48_buf           = pc_w48;


wire                             spc49_inst_done_buf  = spc49_inst_done;
wire [63:0]                      pc_w49_buf           = pc_w49;


wire                             spc50_inst_done_buf  = spc50_inst_done;
wire [63:0]                      pc_w50_buf           = pc_w50;


wire                             spc51_inst_done_buf  = spc51_inst_done;
wire [63:0]                      pc_w51_buf           = pc_w51;


wire                             spc52_inst_done_buf  = spc52_inst_done;
wire [63:0]                      pc_w52_buf           = pc_w52;


wire                             spc53_inst_done_buf  = spc53_inst_done;
wire [63:0]                      pc_w53_buf           = pc_w53;


wire                             spc54_inst_done_buf  = spc54_inst_done;
wire [63:0]                      pc_w54_buf           = pc_w54;


wire                             spc55_inst_done_buf  = spc55_inst_done;
wire [63:0]                      pc_w55_buf           = pc_w55;


wire                             spc56_inst_done_buf  = spc56_inst_done;
wire [63:0]                      pc_w56_buf           = pc_w56;


wire                             spc57_inst_done_buf  = spc57_inst_done;
wire [63:0]                      pc_w57_buf           = pc_w57;


wire                             spc58_inst_done_buf  = spc58_inst_done;
wire [63:0]                      pc_w58_buf           = pc_w58;


wire                             spc59_inst_done_buf  = spc59_inst_done;
wire [63:0]                      pc_w59_buf           = pc_w59;


wire                             spc60_inst_done_buf  = spc60_inst_done;
wire [63:0]                      pc_w60_buf           = pc_w60;


wire                             spc61_inst_done_buf  = spc61_inst_done;
wire [63:0]                      pc_w61_buf           = pc_w61;


wire                             spc62_inst_done_buf  = spc62_inst_done;
wire [63:0]                      pc_w62_buf           = pc_w62;


wire                             spc63_inst_done_buf  = spc63_inst_done;
wire [63:0]                      pc_w63_buf           = pc_w63;


wire                             spc64_inst_done_buf  = spc64_inst_done;
wire [63:0]                      pc_w64_buf           = pc_w64;


wire                             spc65_inst_done_buf  = spc65_inst_done;
wire [63:0]                      pc_w65_buf           = pc_w65;


wire                             spc66_inst_done_buf  = spc66_inst_done;
wire [63:0]                      pc_w66_buf           = pc_w66;


wire                             spc67_inst_done_buf  = spc67_inst_done;
wire [63:0]                      pc_w67_buf           = pc_w67;


wire                             spc68_inst_done_buf  = spc68_inst_done;
wire [63:0]                      pc_w68_buf           = pc_w68;


wire                             spc69_inst_done_buf  = spc69_inst_done;
wire [63:0]                      pc_w69_buf           = pc_w69;


wire                             spc70_inst_done_buf  = spc70_inst_done;
wire [63:0]                      pc_w70_buf           = pc_w70;


wire                             spc71_inst_done_buf  = spc71_inst_done;
wire [63:0]                      pc_w71_buf           = pc_w71;


wire                             spc72_inst_done_buf  = spc72_inst_done;
wire [63:0]                      pc_w72_buf           = pc_w72;


wire                             spc73_inst_done_buf  = spc73_inst_done;
wire [63:0]                      pc_w73_buf           = pc_w73;


wire                             spc74_inst_done_buf  = spc74_inst_done;
wire [63:0]                      pc_w74_buf           = pc_w74;


wire                             spc75_inst_done_buf  = spc75_inst_done;
wire [63:0]                      pc_w75_buf           = pc_w75;


wire                             spc76_inst_done_buf  = spc76_inst_done;
wire [63:0]                      pc_w76_buf           = pc_w76;


wire                             spc77_inst_done_buf  = spc77_inst_done;
wire [63:0]                      pc_w77_buf           = pc_w77;


wire                             spc78_inst_done_buf  = spc78_inst_done;
wire [63:0]                      pc_w78_buf           = pc_w78;


wire                             spc79_inst_done_buf  = spc79_inst_done;
wire [63:0]                      pc_w79_buf           = pc_w79;


wire                             spc80_inst_done_buf  = spc80_inst_done;
wire [63:0]                      pc_w80_buf           = pc_w80;


wire                             spc81_inst_done_buf  = spc81_inst_done;
wire [63:0]                      pc_w81_buf           = pc_w81;


wire                             spc82_inst_done_buf  = spc82_inst_done;
wire [63:0]                      pc_w82_buf           = pc_w82;


wire                             spc83_inst_done_buf  = spc83_inst_done;
wire [63:0]                      pc_w83_buf           = pc_w83;


wire                             spc84_inst_done_buf  = spc84_inst_done;
wire [63:0]                      pc_w84_buf           = pc_w84;


wire                             spc85_inst_done_buf  = spc85_inst_done;
wire [63:0]                      pc_w85_buf           = pc_w85;


wire                             spc86_inst_done_buf  = spc86_inst_done;
wire [63:0]                      pc_w86_buf           = pc_w86;


wire                             spc87_inst_done_buf  = spc87_inst_done;
wire [63:0]                      pc_w87_buf           = pc_w87;


wire                             spc88_inst_done_buf  = spc88_inst_done;
wire [63:0]                      pc_w88_buf           = pc_w88;


wire                             spc89_inst_done_buf  = spc89_inst_done;
wire [63:0]                      pc_w89_buf           = pc_w89;


wire                             spc90_inst_done_buf  = spc90_inst_done;
wire [63:0]                      pc_w90_buf           = pc_w90;


wire                             spc91_inst_done_buf  = spc91_inst_done;
wire [63:0]                      pc_w91_buf           = pc_w91;


wire                             spc92_inst_done_buf  = spc92_inst_done;
wire [63:0]                      pc_w92_buf           = pc_w92;


wire                             spc93_inst_done_buf  = spc93_inst_done;
wire [63:0]                      pc_w93_buf           = pc_w93;


wire                             spc94_inst_done_buf  = spc94_inst_done;
wire [63:0]                      pc_w94_buf           = pc_w94;


wire                             spc95_inst_done_buf  = spc95_inst_done;
wire [63:0]                      pc_w95_buf           = pc_w95;


wire                             spc96_inst_done_buf  = spc96_inst_done;
wire [63:0]                      pc_w96_buf           = pc_w96;


wire                             spc97_inst_done_buf  = spc97_inst_done;
wire [63:0]                      pc_w97_buf           = pc_w97;


wire                             spc98_inst_done_buf  = spc98_inst_done;
wire [63:0]                      pc_w98_buf           = pc_w98;


wire                             spc99_inst_done_buf  = spc99_inst_done;
wire [63:0]                      pc_w99_buf           = pc_w99;


wire                             spc100_inst_done_buf  = spc100_inst_done;
wire [63:0]                      pc_w100_buf           = pc_w100;


wire                             spc101_inst_done_buf  = spc101_inst_done;
wire [63:0]                      pc_w101_buf           = pc_w101;


wire                             spc102_inst_done_buf  = spc102_inst_done;
wire [63:0]                      pc_w102_buf           = pc_w102;


wire                             spc103_inst_done_buf  = spc103_inst_done;
wire [63:0]                      pc_w103_buf           = pc_w103;


wire                             spc104_inst_done_buf  = spc104_inst_done;
wire [63:0]                      pc_w104_buf           = pc_w104;


wire                             spc105_inst_done_buf  = spc105_inst_done;
wire [63:0]                      pc_w105_buf           = pc_w105;


wire                             spc106_inst_done_buf  = spc106_inst_done;
wire [63:0]                      pc_w106_buf           = pc_w106;


wire                             spc107_inst_done_buf  = spc107_inst_done;
wire [63:0]                      pc_w107_buf           = pc_w107;


wire                             spc108_inst_done_buf  = spc108_inst_done;
wire [63:0]                      pc_w108_buf           = pc_w108;


wire                             spc109_inst_done_buf  = spc109_inst_done;
wire [63:0]                      pc_w109_buf           = pc_w109;


wire                             spc110_inst_done_buf  = spc110_inst_done;
wire [63:0]                      pc_w110_buf           = pc_w110;


wire                             spc111_inst_done_buf  = spc111_inst_done;
wire [63:0]                      pc_w111_buf           = pc_w111;


wire                             spc112_inst_done_buf  = spc112_inst_done;
wire [63:0]                      pc_w112_buf           = pc_w112;


wire                             spc113_inst_done_buf  = spc113_inst_done;
wire [63:0]                      pc_w113_buf           = pc_w113;


wire                             spc114_inst_done_buf  = spc114_inst_done;
wire [63:0]                      pc_w114_buf           = pc_w114;


wire                             spc115_inst_done_buf  = spc115_inst_done;
wire [63:0]                      pc_w115_buf           = pc_w115;


wire                             spc116_inst_done_buf  = spc116_inst_done;
wire [63:0]                      pc_w116_buf           = pc_w116;


wire                             spc117_inst_done_buf  = spc117_inst_done;
wire [63:0]                      pc_w117_buf           = pc_w117;


wire                             spc118_inst_done_buf  = spc118_inst_done;
wire [63:0]                      pc_w118_buf           = pc_w118;


wire                             spc119_inst_done_buf  = spc119_inst_done;
wire [63:0]                      pc_w119_buf           = pc_w119;


wire                             spc120_inst_done_buf  = spc120_inst_done;
wire [63:0]                      pc_w120_buf           = pc_w120;


wire                             spc121_inst_done_buf  = spc121_inst_done;
wire [63:0]                      pc_w121_buf           = pc_w121;


wire                             spc122_inst_done_buf  = spc122_inst_done;
wire [63:0]                      pc_w122_buf           = pc_w122;


wire                             spc123_inst_done_buf  = spc123_inst_done;
wire [63:0]                      pc_w123_buf           = pc_w123;


wire                             spc124_inst_done_buf  = spc124_inst_done;
wire [63:0]                      pc_w124_buf           = pc_w124;


wire                             spc125_inst_done_buf  = spc125_inst_done;
wire [63:0]                      pc_w125_buf           = pc_w125;


wire                             spc126_inst_done_buf  = spc126_inst_done;
wire [63:0]                      pc_w126_buf           = pc_w126;


wire                             spc127_inst_done_buf  = spc127_inst_done;
wire [63:0]                      pc_w127_buf           = pc_w127;


wire                             spc128_inst_done_buf  = spc128_inst_done;
wire [63:0]                      pc_w128_buf           = pc_w128;


wire                             spc129_inst_done_buf  = spc129_inst_done;
wire [63:0]                      pc_w129_buf           = pc_w129;


wire                             spc130_inst_done_buf  = spc130_inst_done;
wire [63:0]                      pc_w130_buf           = pc_w130;


wire                             spc131_inst_done_buf  = spc131_inst_done;
wire [63:0]                      pc_w131_buf           = pc_w131;


wire                             spc132_inst_done_buf  = spc132_inst_done;
wire [63:0]                      pc_w132_buf           = pc_w132;


wire                             spc133_inst_done_buf  = spc133_inst_done;
wire [63:0]                      pc_w133_buf           = pc_w133;


wire                             spc134_inst_done_buf  = spc134_inst_done;
wire [63:0]                      pc_w134_buf           = pc_w134;


wire                             spc135_inst_done_buf  = spc135_inst_done;
wire [63:0]                      pc_w135_buf           = pc_w135;


wire                             spc136_inst_done_buf  = spc136_inst_done;
wire [63:0]                      pc_w136_buf           = pc_w136;


wire                             spc137_inst_done_buf  = spc137_inst_done;
wire [63:0]                      pc_w137_buf           = pc_w137;


wire                             spc138_inst_done_buf  = spc138_inst_done;
wire [63:0]                      pc_w138_buf           = pc_w138;


wire                             spc139_inst_done_buf  = spc139_inst_done;
wire [63:0]                      pc_w139_buf           = pc_w139;


wire                             spc140_inst_done_buf  = spc140_inst_done;
wire [63:0]                      pc_w140_buf           = pc_w140;


wire                             spc141_inst_done_buf  = spc141_inst_done;
wire [63:0]                      pc_w141_buf           = pc_w141;


wire                             spc142_inst_done_buf  = spc142_inst_done;
wire [63:0]                      pc_w142_buf           = pc_w142;


wire                             spc143_inst_done_buf  = spc143_inst_done;
wire [63:0]                      pc_w143_buf           = pc_w143;


wire                             spc144_inst_done_buf  = spc144_inst_done;
wire [63:0]                      pc_w144_buf           = pc_w144;


wire                             spc145_inst_done_buf  = spc145_inst_done;
wire [63:0]                      pc_w145_buf           = pc_w145;


wire                             spc146_inst_done_buf  = spc146_inst_done;
wire [63:0]                      pc_w146_buf           = pc_w146;


wire                             spc147_inst_done_buf  = spc147_inst_done;
wire [63:0]                      pc_w147_buf           = pc_w147;


wire                             spc148_inst_done_buf  = spc148_inst_done;
wire [63:0]                      pc_w148_buf           = pc_w148;


wire                             spc149_inst_done_buf  = spc149_inst_done;
wire [63:0]                      pc_w149_buf           = pc_w149;


wire                             spc150_inst_done_buf  = spc150_inst_done;
wire [63:0]                      pc_w150_buf           = pc_w150;


wire                             spc151_inst_done_buf  = spc151_inst_done;
wire [63:0]                      pc_w151_buf           = pc_w151;


wire                             spc152_inst_done_buf  = spc152_inst_done;
wire [63:0]                      pc_w152_buf           = pc_w152;


wire                             spc153_inst_done_buf  = spc153_inst_done;
wire [63:0]                      pc_w153_buf           = pc_w153;


wire                             spc154_inst_done_buf  = spc154_inst_done;
wire [63:0]                      pc_w154_buf           = pc_w154;


wire                             spc155_inst_done_buf  = spc155_inst_done;
wire [63:0]                      pc_w155_buf           = pc_w155;


wire                             spc156_inst_done_buf  = spc156_inst_done;
wire [63:0]                      pc_w156_buf           = pc_w156;


wire                             spc157_inst_done_buf  = spc157_inst_done;
wire [63:0]                      pc_w157_buf           = pc_w157;


wire                             spc158_inst_done_buf  = spc158_inst_done;
wire [63:0]                      pc_w158_buf           = pc_w158;


wire                             spc159_inst_done_buf  = spc159_inst_done;
wire [63:0]                      pc_w159_buf           = pc_w159;


wire                             spc160_inst_done_buf  = spc160_inst_done;
wire [63:0]                      pc_w160_buf           = pc_w160;


wire                             spc161_inst_done_buf  = spc161_inst_done;
wire [63:0]                      pc_w161_buf           = pc_w161;


wire                             spc162_inst_done_buf  = spc162_inst_done;
wire [63:0]                      pc_w162_buf           = pc_w162;


wire                             spc163_inst_done_buf  = spc163_inst_done;
wire [63:0]                      pc_w163_buf           = pc_w163;


wire                             spc164_inst_done_buf  = spc164_inst_done;
wire [63:0]                      pc_w164_buf           = pc_w164;


wire                             spc165_inst_done_buf  = spc165_inst_done;
wire [63:0]                      pc_w165_buf           = pc_w165;


wire                             spc166_inst_done_buf  = spc166_inst_done;
wire [63:0]                      pc_w166_buf           = pc_w166;


wire                             spc167_inst_done_buf  = spc167_inst_done;
wire [63:0]                      pc_w167_buf           = pc_w167;


wire                             spc168_inst_done_buf  = spc168_inst_done;
wire [63:0]                      pc_w168_buf           = pc_w168;


wire                             spc169_inst_done_buf  = spc169_inst_done;
wire [63:0]                      pc_w169_buf           = pc_w169;


wire                             spc170_inst_done_buf  = spc170_inst_done;
wire [63:0]                      pc_w170_buf           = pc_w170;


wire                             spc171_inst_done_buf  = spc171_inst_done;
wire [63:0]                      pc_w171_buf           = pc_w171;


wire                             spc172_inst_done_buf  = spc172_inst_done;
wire [63:0]                      pc_w172_buf           = pc_w172;


wire                             spc173_inst_done_buf  = spc173_inst_done;
wire [63:0]                      pc_w173_buf           = pc_w173;


wire                             spc174_inst_done_buf  = spc174_inst_done;
wire [63:0]                      pc_w174_buf           = pc_w174;


wire                             spc175_inst_done_buf  = spc175_inst_done;
wire [63:0]                      pc_w175_buf           = pc_w175;


wire                             spc176_inst_done_buf  = spc176_inst_done;
wire [63:0]                      pc_w176_buf           = pc_w176;


wire                             spc177_inst_done_buf  = spc177_inst_done;
wire [63:0]                      pc_w177_buf           = pc_w177;


wire                             spc178_inst_done_buf  = spc178_inst_done;
wire [63:0]                      pc_w178_buf           = pc_w178;


wire                             spc179_inst_done_buf  = spc179_inst_done;
wire [63:0]                      pc_w179_buf           = pc_w179;


wire                             spc180_inst_done_buf  = spc180_inst_done;
wire [63:0]                      pc_w180_buf           = pc_w180;


wire                             spc181_inst_done_buf  = spc181_inst_done;
wire [63:0]                      pc_w181_buf           = pc_w181;


wire                             spc182_inst_done_buf  = spc182_inst_done;
wire [63:0]                      pc_w182_buf           = pc_w182;


wire                             spc183_inst_done_buf  = spc183_inst_done;
wire [63:0]                      pc_w183_buf           = pc_w183;


wire                             spc184_inst_done_buf  = spc184_inst_done;
wire [63:0]                      pc_w184_buf           = pc_w184;


wire                             spc185_inst_done_buf  = spc185_inst_done;
wire [63:0]                      pc_w185_buf           = pc_w185;


wire                             spc186_inst_done_buf  = spc186_inst_done;
wire [63:0]                      pc_w186_buf           = pc_w186;


wire                             spc187_inst_done_buf  = spc187_inst_done;
wire [63:0]                      pc_w187_buf           = pc_w187;


wire                             spc188_inst_done_buf  = spc188_inst_done;
wire [63:0]                      pc_w188_buf           = pc_w188;


wire                             spc189_inst_done_buf  = spc189_inst_done;
wire [63:0]                      pc_w189_buf           = pc_w189;


wire                             spc190_inst_done_buf  = spc190_inst_done;
wire [63:0]                      pc_w190_buf           = pc_w190;


wire                             spc191_inst_done_buf  = spc191_inst_done;
wire [63:0]                      pc_w191_buf           = pc_w191;


wire                             spc192_inst_done_buf  = spc192_inst_done;
wire [63:0]                      pc_w192_buf           = pc_w192;


wire                             spc193_inst_done_buf  = spc193_inst_done;
wire [63:0]                      pc_w193_buf           = pc_w193;


wire                             spc194_inst_done_buf  = spc194_inst_done;
wire [63:0]                      pc_w194_buf           = pc_w194;


wire                             spc195_inst_done_buf  = spc195_inst_done;
wire [63:0]                      pc_w195_buf           = pc_w195;


wire                             spc196_inst_done_buf  = spc196_inst_done;
wire [63:0]                      pc_w196_buf           = pc_w196;


wire                             spc197_inst_done_buf  = spc197_inst_done;
wire [63:0]                      pc_w197_buf           = pc_w197;


wire                             spc198_inst_done_buf  = spc198_inst_done;
wire [63:0]                      pc_w198_buf           = pc_w198;


wire                             spc199_inst_done_buf  = spc199_inst_done;
wire [63:0]                      pc_w199_buf           = pc_w199;


wire                             spc200_inst_done_buf  = spc200_inst_done;
wire [63:0]                      pc_w200_buf           = pc_w200;


wire                             spc201_inst_done_buf  = spc201_inst_done;
wire [63:0]                      pc_w201_buf           = pc_w201;


wire                             spc202_inst_done_buf  = spc202_inst_done;
wire [63:0]                      pc_w202_buf           = pc_w202;


wire                             spc203_inst_done_buf  = spc203_inst_done;
wire [63:0]                      pc_w203_buf           = pc_w203;


wire                             spc204_inst_done_buf  = spc204_inst_done;
wire [63:0]                      pc_w204_buf           = pc_w204;


wire                             spc205_inst_done_buf  = spc205_inst_done;
wire [63:0]                      pc_w205_buf           = pc_w205;


wire                             spc206_inst_done_buf  = spc206_inst_done;
wire [63:0]                      pc_w206_buf           = pc_w206;


wire                             spc207_inst_done_buf  = spc207_inst_done;
wire [63:0]                      pc_w207_buf           = pc_w207;


wire                             spc208_inst_done_buf  = spc208_inst_done;
wire [63:0]                      pc_w208_buf           = pc_w208;


wire                             spc209_inst_done_buf  = spc209_inst_done;
wire [63:0]                      pc_w209_buf           = pc_w209;


wire                             spc210_inst_done_buf  = spc210_inst_done;
wire [63:0]                      pc_w210_buf           = pc_w210;


wire                             spc211_inst_done_buf  = spc211_inst_done;
wire [63:0]                      pc_w211_buf           = pc_w211;


wire                             spc212_inst_done_buf  = spc212_inst_done;
wire [63:0]                      pc_w212_buf           = pc_w212;


wire                             spc213_inst_done_buf  = spc213_inst_done;
wire [63:0]                      pc_w213_buf           = pc_w213;


wire                             spc214_inst_done_buf  = spc214_inst_done;
wire [63:0]                      pc_w214_buf           = pc_w214;


wire                             spc215_inst_done_buf  = spc215_inst_done;
wire [63:0]                      pc_w215_buf           = pc_w215;


wire                             spc216_inst_done_buf  = spc216_inst_done;
wire [63:0]                      pc_w216_buf           = pc_w216;


wire                             spc217_inst_done_buf  = spc217_inst_done;
wire [63:0]                      pc_w217_buf           = pc_w217;


wire                             spc218_inst_done_buf  = spc218_inst_done;
wire [63:0]                      pc_w218_buf           = pc_w218;


wire                             spc219_inst_done_buf  = spc219_inst_done;
wire [63:0]                      pc_w219_buf           = pc_w219;


wire                             spc220_inst_done_buf  = spc220_inst_done;
wire [63:0]                      pc_w220_buf           = pc_w220;


wire                             spc221_inst_done_buf  = spc221_inst_done;
wire [63:0]                      pc_w221_buf           = pc_w221;


wire                             spc222_inst_done_buf  = spc222_inst_done;
wire [63:0]                      pc_w222_buf           = pc_w222;


wire                             spc223_inst_done_buf  = spc223_inst_done;
wire [63:0]                      pc_w223_buf           = pc_w223;


wire                             spc224_inst_done_buf  = spc224_inst_done;
wire [63:0]                      pc_w224_buf           = pc_w224;


wire                             spc225_inst_done_buf  = spc225_inst_done;
wire [63:0]                      pc_w225_buf           = pc_w225;


wire                             spc226_inst_done_buf  = spc226_inst_done;
wire [63:0]                      pc_w226_buf           = pc_w226;


wire                             spc227_inst_done_buf  = spc227_inst_done;
wire [63:0]                      pc_w227_buf           = pc_w227;


wire                             spc228_inst_done_buf  = spc228_inst_done;
wire [63:0]                      pc_w228_buf           = pc_w228;


wire                             spc229_inst_done_buf  = spc229_inst_done;
wire [63:0]                      pc_w229_buf           = pc_w229;


wire                             spc230_inst_done_buf  = spc230_inst_done;
wire [63:0]                      pc_w230_buf           = pc_w230;


wire                             spc231_inst_done_buf  = spc231_inst_done;
wire [63:0]                      pc_w231_buf           = pc_w231;


wire                             spc232_inst_done_buf  = spc232_inst_done;
wire [63:0]                      pc_w232_buf           = pc_w232;


wire                             spc233_inst_done_buf  = spc233_inst_done;
wire [63:0]                      pc_w233_buf           = pc_w233;


wire                             spc234_inst_done_buf  = spc234_inst_done;
wire [63:0]                      pc_w234_buf           = pc_w234;


wire                             spc235_inst_done_buf  = spc235_inst_done;
wire [63:0]                      pc_w235_buf           = pc_w235;


wire                             spc236_inst_done_buf  = spc236_inst_done;
wire [63:0]                      pc_w236_buf           = pc_w236;


wire                             spc237_inst_done_buf  = spc237_inst_done;
wire [63:0]                      pc_w237_buf           = pc_w237;


wire                             spc238_inst_done_buf  = spc238_inst_done;
wire [63:0]                      pc_w238_buf           = pc_w238;


wire                             spc239_inst_done_buf  = spc239_inst_done;
wire [63:0]                      pc_w239_buf           = pc_w239;


wire                             spc240_inst_done_buf  = spc240_inst_done;
wire [63:0]                      pc_w240_buf           = pc_w240;


wire                             spc241_inst_done_buf  = spc241_inst_done;
wire [63:0]                      pc_w241_buf           = pc_w241;


wire                             spc242_inst_done_buf  = spc242_inst_done;
wire [63:0]                      pc_w242_buf           = pc_w242;


wire                             spc243_inst_done_buf  = spc243_inst_done;
wire [63:0]                      pc_w243_buf           = pc_w243;


wire                             spc244_inst_done_buf  = spc244_inst_done;
wire [63:0]                      pc_w244_buf           = pc_w244;


wire                             spc245_inst_done_buf  = spc245_inst_done;
wire [63:0]                      pc_w245_buf           = pc_w245;


wire                             spc246_inst_done_buf  = spc246_inst_done;
wire [63:0]                      pc_w246_buf           = pc_w246;


wire                             spc247_inst_done_buf  = spc247_inst_done;
wire [63:0]                      pc_w247_buf           = pc_w247;


wire                             spc248_inst_done_buf  = spc248_inst_done;
wire [63:0]                      pc_w248_buf           = pc_w248;


wire                             spc249_inst_done_buf  = spc249_inst_done;
wire [63:0]                      pc_w249_buf           = pc_w249;


wire                             spc250_inst_done_buf  = spc250_inst_done;
wire [63:0]                      pc_w250_buf           = pc_w250;


wire                             spc251_inst_done_buf  = spc251_inst_done;
wire [63:0]                      pc_w251_buf           = pc_w251;


wire                             spc252_inst_done_buf  = spc252_inst_done;
wire [63:0]                      pc_w252_buf           = pc_w252;


wire                             spc253_inst_done_buf  = spc253_inst_done;
wire [63:0]                      pc_w253_buf           = pc_w253;


wire                             spc254_inst_done_buf  = spc254_inst_done;
wire [63:0]                      pc_w254_buf           = pc_w254;


wire                             spc255_inst_done_buf  = spc255_inst_done;
wire [63:0]                      pc_w255_buf           = pc_w255;


wire                             spc256_inst_done_buf  = spc256_inst_done;
wire [63:0]                      pc_w256_buf           = pc_w256;


wire                             spc257_inst_done_buf  = spc257_inst_done;
wire [63:0]                      pc_w257_buf           = pc_w257;


wire                             spc258_inst_done_buf  = spc258_inst_done;
wire [63:0]                      pc_w258_buf           = pc_w258;


wire                             spc259_inst_done_buf  = spc259_inst_done;
wire [63:0]                      pc_w259_buf           = pc_w259;


wire                             spc260_inst_done_buf  = spc260_inst_done;
wire [63:0]                      pc_w260_buf           = pc_w260;


wire                             spc261_inst_done_buf  = spc261_inst_done;
wire [63:0]                      pc_w261_buf           = pc_w261;


wire                             spc262_inst_done_buf  = spc262_inst_done;
wire [63:0]                      pc_w262_buf           = pc_w262;


wire                             spc263_inst_done_buf  = spc263_inst_done;
wire [63:0]                      pc_w263_buf           = pc_w263;


wire                             spc264_inst_done_buf  = spc264_inst_done;
wire [63:0]                      pc_w264_buf           = pc_w264;


wire                             spc265_inst_done_buf  = spc265_inst_done;
wire [63:0]                      pc_w265_buf           = pc_w265;


wire                             spc266_inst_done_buf  = spc266_inst_done;
wire [63:0]                      pc_w266_buf           = pc_w266;


wire                             spc267_inst_done_buf  = spc267_inst_done;
wire [63:0]                      pc_w267_buf           = pc_w267;


wire                             spc268_inst_done_buf  = spc268_inst_done;
wire [63:0]                      pc_w268_buf           = pc_w268;


wire                             spc269_inst_done_buf  = spc269_inst_done;
wire [63:0]                      pc_w269_buf           = pc_w269;


wire                             spc270_inst_done_buf  = spc270_inst_done;
wire [63:0]                      pc_w270_buf           = pc_w270;


wire                             spc271_inst_done_buf  = spc271_inst_done;
wire [63:0]                      pc_w271_buf           = pc_w271;


wire                             spc272_inst_done_buf  = spc272_inst_done;
wire [63:0]                      pc_w272_buf           = pc_w272;


wire                             spc273_inst_done_buf  = spc273_inst_done;
wire [63:0]                      pc_w273_buf           = pc_w273;


wire                             spc274_inst_done_buf  = spc274_inst_done;
wire [63:0]                      pc_w274_buf           = pc_w274;


wire                             spc275_inst_done_buf  = spc275_inst_done;
wire [63:0]                      pc_w275_buf           = pc_w275;


wire                             spc276_inst_done_buf  = spc276_inst_done;
wire [63:0]                      pc_w276_buf           = pc_w276;


wire                             spc277_inst_done_buf  = spc277_inst_done;
wire [63:0]                      pc_w277_buf           = pc_w277;


wire                             spc278_inst_done_buf  = spc278_inst_done;
wire [63:0]                      pc_w278_buf           = pc_w278;


wire                             spc279_inst_done_buf  = spc279_inst_done;
wire [63:0]                      pc_w279_buf           = pc_w279;


wire                             spc280_inst_done_buf  = spc280_inst_done;
wire [63:0]                      pc_w280_buf           = pc_w280;


wire                             spc281_inst_done_buf  = spc281_inst_done;
wire [63:0]                      pc_w281_buf           = pc_w281;


wire                             spc282_inst_done_buf  = spc282_inst_done;
wire [63:0]                      pc_w282_buf           = pc_w282;


wire                             spc283_inst_done_buf  = spc283_inst_done;
wire [63:0]                      pc_w283_buf           = pc_w283;


wire                             spc284_inst_done_buf  = spc284_inst_done;
wire [63:0]                      pc_w284_buf           = pc_w284;


wire                             spc285_inst_done_buf  = spc285_inst_done;
wire [63:0]                      pc_w285_buf           = pc_w285;


wire                             spc286_inst_done_buf  = spc286_inst_done;
wire [63:0]                      pc_w286_buf           = pc_w286;


wire                             spc287_inst_done_buf  = spc287_inst_done;
wire [63:0]                      pc_w287_buf           = pc_w287;


wire                             spc288_inst_done_buf  = spc288_inst_done;
wire [63:0]                      pc_w288_buf           = pc_w288;


wire                             spc289_inst_done_buf  = spc289_inst_done;
wire [63:0]                      pc_w289_buf           = pc_w289;


wire                             spc290_inst_done_buf  = spc290_inst_done;
wire [63:0]                      pc_w290_buf           = pc_w290;


wire                             spc291_inst_done_buf  = spc291_inst_done;
wire [63:0]                      pc_w291_buf           = pc_w291;


wire                             spc292_inst_done_buf  = spc292_inst_done;
wire [63:0]                      pc_w292_buf           = pc_w292;


wire                             spc293_inst_done_buf  = spc293_inst_done;
wire [63:0]                      pc_w293_buf           = pc_w293;


wire                             spc294_inst_done_buf  = spc294_inst_done;
wire [63:0]                      pc_w294_buf           = pc_w294;


wire                             spc295_inst_done_buf  = spc295_inst_done;
wire [63:0]                      pc_w295_buf           = pc_w295;


wire                             spc296_inst_done_buf  = spc296_inst_done;
wire [63:0]                      pc_w296_buf           = pc_w296;


wire                             spc297_inst_done_buf  = spc297_inst_done;
wire [63:0]                      pc_w297_buf           = pc_w297;


wire                             spc298_inst_done_buf  = spc298_inst_done;
wire [63:0]                      pc_w298_buf           = pc_w298;


wire                             spc299_inst_done_buf  = spc299_inst_done;
wire [63:0]                      pc_w299_buf           = pc_w299;


wire                             spc300_inst_done_buf  = spc300_inst_done;
wire [63:0]                      pc_w300_buf           = pc_w300;


wire                             spc301_inst_done_buf  = spc301_inst_done;
wire [63:0]                      pc_w301_buf           = pc_w301;


wire                             spc302_inst_done_buf  = spc302_inst_done;
wire [63:0]                      pc_w302_buf           = pc_w302;


wire                             spc303_inst_done_buf  = spc303_inst_done;
wire [63:0]                      pc_w303_buf           = pc_w303;


wire                             spc304_inst_done_buf  = spc304_inst_done;
wire [63:0]                      pc_w304_buf           = pc_w304;


wire                             spc305_inst_done_buf  = spc305_inst_done;
wire [63:0]                      pc_w305_buf           = pc_w305;


wire                             spc306_inst_done_buf  = spc306_inst_done;
wire [63:0]                      pc_w306_buf           = pc_w306;


wire                             spc307_inst_done_buf  = spc307_inst_done;
wire [63:0]                      pc_w307_buf           = pc_w307;


wire                             spc308_inst_done_buf  = spc308_inst_done;
wire [63:0]                      pc_w308_buf           = pc_w308;


wire                             spc309_inst_done_buf  = spc309_inst_done;
wire [63:0]                      pc_w309_buf           = pc_w309;


wire                             spc310_inst_done_buf  = spc310_inst_done;
wire [63:0]                      pc_w310_buf           = pc_w310;


wire                             spc311_inst_done_buf  = spc311_inst_done;
wire [63:0]                      pc_w311_buf           = pc_w311;


wire                             spc312_inst_done_buf  = spc312_inst_done;
wire [63:0]                      pc_w312_buf           = pc_w312;


wire                             spc313_inst_done_buf  = spc313_inst_done;
wire [63:0]                      pc_w313_buf           = pc_w313;


wire                             spc314_inst_done_buf  = spc314_inst_done;
wire [63:0]                      pc_w314_buf           = pc_w314;


wire                             spc315_inst_done_buf  = spc315_inst_done;
wire [63:0]                      pc_w315_buf           = pc_w315;


wire                             spc316_inst_done_buf  = spc316_inst_done;
wire [63:0]                      pc_w316_buf           = pc_w316;


wire                             spc317_inst_done_buf  = spc317_inst_done;
wire [63:0]                      pc_w317_buf           = pc_w317;


wire                             spc318_inst_done_buf  = spc318_inst_done;
wire [63:0]                      pc_w318_buf           = pc_w318;


wire                             spc319_inst_done_buf  = spc319_inst_done;
wire [63:0]                      pc_w319_buf           = pc_w319;


wire                             spc320_inst_done_buf  = spc320_inst_done;
wire [63:0]                      pc_w320_buf           = pc_w320;


wire                             spc321_inst_done_buf  = spc321_inst_done;
wire [63:0]                      pc_w321_buf           = pc_w321;


wire                             spc322_inst_done_buf  = spc322_inst_done;
wire [63:0]                      pc_w322_buf           = pc_w322;


wire                             spc323_inst_done_buf  = spc323_inst_done;
wire [63:0]                      pc_w323_buf           = pc_w323;


wire                             spc324_inst_done_buf  = spc324_inst_done;
wire [63:0]                      pc_w324_buf           = pc_w324;


wire                             spc325_inst_done_buf  = spc325_inst_done;
wire [63:0]                      pc_w325_buf           = pc_w325;


wire                             spc326_inst_done_buf  = spc326_inst_done;
wire [63:0]                      pc_w326_buf           = pc_w326;


wire                             spc327_inst_done_buf  = spc327_inst_done;
wire [63:0]                      pc_w327_buf           = pc_w327;


wire                             spc328_inst_done_buf  = spc328_inst_done;
wire [63:0]                      pc_w328_buf           = pc_w328;


wire                             spc329_inst_done_buf  = spc329_inst_done;
wire [63:0]                      pc_w329_buf           = pc_w329;


wire                             spc330_inst_done_buf  = spc330_inst_done;
wire [63:0]                      pc_w330_buf           = pc_w330;


wire                             spc331_inst_done_buf  = spc331_inst_done;
wire [63:0]                      pc_w331_buf           = pc_w331;


wire                             spc332_inst_done_buf  = spc332_inst_done;
wire [63:0]                      pc_w332_buf           = pc_w332;


wire                             spc333_inst_done_buf  = spc333_inst_done;
wire [63:0]                      pc_w333_buf           = pc_w333;


wire                             spc334_inst_done_buf  = spc334_inst_done;
wire [63:0]                      pc_w334_buf           = pc_w334;


wire                             spc335_inst_done_buf  = spc335_inst_done;
wire [63:0]                      pc_w335_buf           = pc_w335;


wire                             spc336_inst_done_buf  = spc336_inst_done;
wire [63:0]                      pc_w336_buf           = pc_w336;


wire                             spc337_inst_done_buf  = spc337_inst_done;
wire [63:0]                      pc_w337_buf           = pc_w337;


wire                             spc338_inst_done_buf  = spc338_inst_done;
wire [63:0]                      pc_w338_buf           = pc_w338;


wire                             spc339_inst_done_buf  = spc339_inst_done;
wire [63:0]                      pc_w339_buf           = pc_w339;


wire                             spc340_inst_done_buf  = spc340_inst_done;
wire [63:0]                      pc_w340_buf           = pc_w340;


wire                             spc341_inst_done_buf  = spc341_inst_done;
wire [63:0]                      pc_w341_buf           = pc_w341;


wire                             spc342_inst_done_buf  = spc342_inst_done;
wire [63:0]                      pc_w342_buf           = pc_w342;


wire                             spc343_inst_done_buf  = spc343_inst_done;
wire [63:0]                      pc_w343_buf           = pc_w343;


wire                             spc344_inst_done_buf  = spc344_inst_done;
wire [63:0]                      pc_w344_buf           = pc_w344;


wire                             spc345_inst_done_buf  = spc345_inst_done;
wire [63:0]                      pc_w345_buf           = pc_w345;


wire                             spc346_inst_done_buf  = spc346_inst_done;
wire [63:0]                      pc_w346_buf           = pc_w346;


wire                             spc347_inst_done_buf  = spc347_inst_done;
wire [63:0]                      pc_w347_buf           = pc_w347;


wire                             spc348_inst_done_buf  = spc348_inst_done;
wire [63:0]                      pc_w348_buf           = pc_w348;


wire                             spc349_inst_done_buf  = spc349_inst_done;
wire [63:0]                      pc_w349_buf           = pc_w349;


wire                             spc350_inst_done_buf  = spc350_inst_done;
wire [63:0]                      pc_w350_buf           = pc_w350;


wire                             spc351_inst_done_buf  = spc351_inst_done;
wire [63:0]                      pc_w351_buf           = pc_w351;


wire                             spc352_inst_done_buf  = spc352_inst_done;
wire [63:0]                      pc_w352_buf           = pc_w352;


wire                             spc353_inst_done_buf  = spc353_inst_done;
wire [63:0]                      pc_w353_buf           = pc_w353;


wire                             spc354_inst_done_buf  = spc354_inst_done;
wire [63:0]                      pc_w354_buf           = pc_w354;


wire                             spc355_inst_done_buf  = spc355_inst_done;
wire [63:0]                      pc_w355_buf           = pc_w355;


wire                             spc356_inst_done_buf  = spc356_inst_done;
wire [63:0]                      pc_w356_buf           = pc_w356;


wire                             spc357_inst_done_buf  = spc357_inst_done;
wire [63:0]                      pc_w357_buf           = pc_w357;


wire                             spc358_inst_done_buf  = spc358_inst_done;
wire [63:0]                      pc_w358_buf           = pc_w358;


wire                             spc359_inst_done_buf  = spc359_inst_done;
wire [63:0]                      pc_w359_buf           = pc_w359;


wire                             spc360_inst_done_buf  = spc360_inst_done;
wire [63:0]                      pc_w360_buf           = pc_w360;


wire                             spc361_inst_done_buf  = spc361_inst_done;
wire [63:0]                      pc_w361_buf           = pc_w361;


wire                             spc362_inst_done_buf  = spc362_inst_done;
wire [63:0]                      pc_w362_buf           = pc_w362;


wire                             spc363_inst_done_buf  = spc363_inst_done;
wire [63:0]                      pc_w363_buf           = pc_w363;


wire                             spc364_inst_done_buf  = spc364_inst_done;
wire [63:0]                      pc_w364_buf           = pc_w364;


wire                             spc365_inst_done_buf  = spc365_inst_done;
wire [63:0]                      pc_w365_buf           = pc_w365;


wire                             spc366_inst_done_buf  = spc366_inst_done;
wire [63:0]                      pc_w366_buf           = pc_w366;


wire                             spc367_inst_done_buf  = spc367_inst_done;
wire [63:0]                      pc_w367_buf           = pc_w367;


wire                             spc368_inst_done_buf  = spc368_inst_done;
wire [63:0]                      pc_w368_buf           = pc_w368;


wire                             spc369_inst_done_buf  = spc369_inst_done;
wire [63:0]                      pc_w369_buf           = pc_w369;


wire                             spc370_inst_done_buf  = spc370_inst_done;
wire [63:0]                      pc_w370_buf           = pc_w370;


wire                             spc371_inst_done_buf  = spc371_inst_done;
wire [63:0]                      pc_w371_buf           = pc_w371;


wire                             spc372_inst_done_buf  = spc372_inst_done;
wire [63:0]                      pc_w372_buf           = pc_w372;


wire                             spc373_inst_done_buf  = spc373_inst_done;
wire [63:0]                      pc_w373_buf           = pc_w373;


wire                             spc374_inst_done_buf  = spc374_inst_done;
wire [63:0]                      pc_w374_buf           = pc_w374;


wire                             spc375_inst_done_buf  = spc375_inst_done;
wire [63:0]                      pc_w375_buf           = pc_w375;


wire                             spc376_inst_done_buf  = spc376_inst_done;
wire [63:0]                      pc_w376_buf           = pc_w376;


wire                             spc377_inst_done_buf  = spc377_inst_done;
wire [63:0]                      pc_w377_buf           = pc_w377;


wire                             spc378_inst_done_buf  = spc378_inst_done;
wire [63:0]                      pc_w378_buf           = pc_w378;


wire                             spc379_inst_done_buf  = spc379_inst_done;
wire [63:0]                      pc_w379_buf           = pc_w379;


wire                             spc380_inst_done_buf  = spc380_inst_done;
wire [63:0]                      pc_w380_buf           = pc_w380;


wire                             spc381_inst_done_buf  = spc381_inst_done;
wire [63:0]                      pc_w381_buf           = pc_w381;


wire                             spc382_inst_done_buf  = spc382_inst_done;
wire [63:0]                      pc_w382_buf           = pc_w382;


wire                             spc383_inst_done_buf  = spc383_inst_done;
wire [63:0]                      pc_w383_buf           = pc_w383;


wire                             spc384_inst_done_buf  = spc384_inst_done;
wire [63:0]                      pc_w384_buf           = pc_w384;


wire                             spc385_inst_done_buf  = spc385_inst_done;
wire [63:0]                      pc_w385_buf           = pc_w385;


wire                             spc386_inst_done_buf  = spc386_inst_done;
wire [63:0]                      pc_w386_buf           = pc_w386;


wire                             spc387_inst_done_buf  = spc387_inst_done;
wire [63:0]                      pc_w387_buf           = pc_w387;


wire                             spc388_inst_done_buf  = spc388_inst_done;
wire [63:0]                      pc_w388_buf           = pc_w388;


wire                             spc389_inst_done_buf  = spc389_inst_done;
wire [63:0]                      pc_w389_buf           = pc_w389;


wire                             spc390_inst_done_buf  = spc390_inst_done;
wire [63:0]                      pc_w390_buf           = pc_w390;


wire                             spc391_inst_done_buf  = spc391_inst_done;
wire [63:0]                      pc_w391_buf           = pc_w391;


wire                             spc392_inst_done_buf  = spc392_inst_done;
wire [63:0]                      pc_w392_buf           = pc_w392;


wire                             spc393_inst_done_buf  = spc393_inst_done;
wire [63:0]                      pc_w393_buf           = pc_w393;


wire                             spc394_inst_done_buf  = spc394_inst_done;
wire [63:0]                      pc_w394_buf           = pc_w394;


wire                             spc395_inst_done_buf  = spc395_inst_done;
wire [63:0]                      pc_w395_buf           = pc_w395;


wire                             spc396_inst_done_buf  = spc396_inst_done;
wire [63:0]                      pc_w396_buf           = pc_w396;


wire                             spc397_inst_done_buf  = spc397_inst_done;
wire [63:0]                      pc_w397_buf           = pc_w397;


wire                             spc398_inst_done_buf  = spc398_inst_done;
wire [63:0]                      pc_w398_buf           = pc_w398;


wire                             spc399_inst_done_buf  = spc399_inst_done;
wire [63:0]                      pc_w399_buf           = pc_w399;


wire                             spc400_inst_done_buf  = spc400_inst_done;
wire [63:0]                      pc_w400_buf           = pc_w400;


wire                             spc401_inst_done_buf  = spc401_inst_done;
wire [63:0]                      pc_w401_buf           = pc_w401;


wire                             spc402_inst_done_buf  = spc402_inst_done;
wire [63:0]                      pc_w402_buf           = pc_w402;


wire                             spc403_inst_done_buf  = spc403_inst_done;
wire [63:0]                      pc_w403_buf           = pc_w403;


wire                             spc404_inst_done_buf  = spc404_inst_done;
wire [63:0]                      pc_w404_buf           = pc_w404;


wire                             spc405_inst_done_buf  = spc405_inst_done;
wire [63:0]                      pc_w405_buf           = pc_w405;


wire                             spc406_inst_done_buf  = spc406_inst_done;
wire [63:0]                      pc_w406_buf           = pc_w406;


wire                             spc407_inst_done_buf  = spc407_inst_done;
wire [63:0]                      pc_w407_buf           = pc_w407;


wire                             spc408_inst_done_buf  = spc408_inst_done;
wire [63:0]                      pc_w408_buf           = pc_w408;


wire                             spc409_inst_done_buf  = spc409_inst_done;
wire [63:0]                      pc_w409_buf           = pc_w409;


wire                             spc410_inst_done_buf  = spc410_inst_done;
wire [63:0]                      pc_w410_buf           = pc_w410;


wire                             spc411_inst_done_buf  = spc411_inst_done;
wire [63:0]                      pc_w411_buf           = pc_w411;


wire                             spc412_inst_done_buf  = spc412_inst_done;
wire [63:0]                      pc_w412_buf           = pc_w412;


wire                             spc413_inst_done_buf  = spc413_inst_done;
wire [63:0]                      pc_w413_buf           = pc_w413;


wire                             spc414_inst_done_buf  = spc414_inst_done;
wire [63:0]                      pc_w414_buf           = pc_w414;


wire                             spc415_inst_done_buf  = spc415_inst_done;
wire [63:0]                      pc_w415_buf           = pc_w415;


wire                             spc416_inst_done_buf  = spc416_inst_done;
wire [63:0]                      pc_w416_buf           = pc_w416;


wire                             spc417_inst_done_buf  = spc417_inst_done;
wire [63:0]                      pc_w417_buf           = pc_w417;


wire                             spc418_inst_done_buf  = spc418_inst_done;
wire [63:0]                      pc_w418_buf           = pc_w418;


wire                             spc419_inst_done_buf  = spc419_inst_done;
wire [63:0]                      pc_w419_buf           = pc_w419;


wire                             spc420_inst_done_buf  = spc420_inst_done;
wire [63:0]                      pc_w420_buf           = pc_w420;


wire                             spc421_inst_done_buf  = spc421_inst_done;
wire [63:0]                      pc_w421_buf           = pc_w421;


wire                             spc422_inst_done_buf  = spc422_inst_done;
wire [63:0]                      pc_w422_buf           = pc_w422;


wire                             spc423_inst_done_buf  = spc423_inst_done;
wire [63:0]                      pc_w423_buf           = pc_w423;


wire                             spc424_inst_done_buf  = spc424_inst_done;
wire [63:0]                      pc_w424_buf           = pc_w424;


wire                             spc425_inst_done_buf  = spc425_inst_done;
wire [63:0]                      pc_w425_buf           = pc_w425;


wire                             spc426_inst_done_buf  = spc426_inst_done;
wire [63:0]                      pc_w426_buf           = pc_w426;


wire                             spc427_inst_done_buf  = spc427_inst_done;
wire [63:0]                      pc_w427_buf           = pc_w427;


wire                             spc428_inst_done_buf  = spc428_inst_done;
wire [63:0]                      pc_w428_buf           = pc_w428;


wire                             spc429_inst_done_buf  = spc429_inst_done;
wire [63:0]                      pc_w429_buf           = pc_w429;


wire                             spc430_inst_done_buf  = spc430_inst_done;
wire [63:0]                      pc_w430_buf           = pc_w430;


wire                             spc431_inst_done_buf  = spc431_inst_done;
wire [63:0]                      pc_w431_buf           = pc_w431;


wire                             spc432_inst_done_buf  = spc432_inst_done;
wire [63:0]                      pc_w432_buf           = pc_w432;


wire                             spc433_inst_done_buf  = spc433_inst_done;
wire [63:0]                      pc_w433_buf           = pc_w433;


wire                             spc434_inst_done_buf  = spc434_inst_done;
wire [63:0]                      pc_w434_buf           = pc_w434;


wire                             spc435_inst_done_buf  = spc435_inst_done;
wire [63:0]                      pc_w435_buf           = pc_w435;


wire                             spc436_inst_done_buf  = spc436_inst_done;
wire [63:0]                      pc_w436_buf           = pc_w436;


wire                             spc437_inst_done_buf  = spc437_inst_done;
wire [63:0]                      pc_w437_buf           = pc_w437;


wire                             spc438_inst_done_buf  = spc438_inst_done;
wire [63:0]                      pc_w438_buf           = pc_w438;


wire                             spc439_inst_done_buf  = spc439_inst_done;
wire [63:0]                      pc_w439_buf           = pc_w439;


wire                             spc440_inst_done_buf  = spc440_inst_done;
wire [63:0]                      pc_w440_buf           = pc_w440;


wire                             spc441_inst_done_buf  = spc441_inst_done;
wire [63:0]                      pc_w441_buf           = pc_w441;


wire                             spc442_inst_done_buf  = spc442_inst_done;
wire [63:0]                      pc_w442_buf           = pc_w442;


wire                             spc443_inst_done_buf  = spc443_inst_done;
wire [63:0]                      pc_w443_buf           = pc_w443;


wire                             spc444_inst_done_buf  = spc444_inst_done;
wire [63:0]                      pc_w444_buf           = pc_w444;


wire                             spc445_inst_done_buf  = spc445_inst_done;
wire [63:0]                      pc_w445_buf           = pc_w445;


wire                             spc446_inst_done_buf  = spc446_inst_done;
wire [63:0]                      pc_w446_buf           = pc_w446;


wire                             spc447_inst_done_buf  = spc447_inst_done;
wire [63:0]                      pc_w447_buf           = pc_w447;


wire                             spc448_inst_done_buf  = spc448_inst_done;
wire [63:0]                      pc_w448_buf           = pc_w448;


wire                             spc449_inst_done_buf  = spc449_inst_done;
wire [63:0]                      pc_w449_buf           = pc_w449;


wire                             spc450_inst_done_buf  = spc450_inst_done;
wire [63:0]                      pc_w450_buf           = pc_w450;


wire                             spc451_inst_done_buf  = spc451_inst_done;
wire [63:0]                      pc_w451_buf           = pc_w451;


wire                             spc452_inst_done_buf  = spc452_inst_done;
wire [63:0]                      pc_w452_buf           = pc_w452;


wire                             spc453_inst_done_buf  = spc453_inst_done;
wire [63:0]                      pc_w453_buf           = pc_w453;


wire                             spc454_inst_done_buf  = spc454_inst_done;
wire [63:0]                      pc_w454_buf           = pc_w454;


wire                             spc455_inst_done_buf  = spc455_inst_done;
wire [63:0]                      pc_w455_buf           = pc_w455;


wire                             spc456_inst_done_buf  = spc456_inst_done;
wire [63:0]                      pc_w456_buf           = pc_w456;


wire                             spc457_inst_done_buf  = spc457_inst_done;
wire [63:0]                      pc_w457_buf           = pc_w457;


wire                             spc458_inst_done_buf  = spc458_inst_done;
wire [63:0]                      pc_w458_buf           = pc_w458;


wire                             spc459_inst_done_buf  = spc459_inst_done;
wire [63:0]                      pc_w459_buf           = pc_w459;


wire                             spc460_inst_done_buf  = spc460_inst_done;
wire [63:0]                      pc_w460_buf           = pc_w460;


wire                             spc461_inst_done_buf  = spc461_inst_done;
wire [63:0]                      pc_w461_buf           = pc_w461;


wire                             spc462_inst_done_buf  = spc462_inst_done;
wire [63:0]                      pc_w462_buf           = pc_w462;


wire                             spc463_inst_done_buf  = spc463_inst_done;
wire [63:0]                      pc_w463_buf           = pc_w463;


wire                             spc464_inst_done_buf  = spc464_inst_done;
wire [63:0]                      pc_w464_buf           = pc_w464;


wire                             spc465_inst_done_buf  = spc465_inst_done;
wire [63:0]                      pc_w465_buf           = pc_w465;


wire                             spc466_inst_done_buf  = spc466_inst_done;
wire [63:0]                      pc_w466_buf           = pc_w466;


wire                             spc467_inst_done_buf  = spc467_inst_done;
wire [63:0]                      pc_w467_buf           = pc_w467;


wire                             spc468_inst_done_buf  = spc468_inst_done;
wire [63:0]                      pc_w468_buf           = pc_w468;


wire                             spc469_inst_done_buf  = spc469_inst_done;
wire [63:0]                      pc_w469_buf           = pc_w469;


wire                             spc470_inst_done_buf  = spc470_inst_done;
wire [63:0]                      pc_w470_buf           = pc_w470;


wire                             spc471_inst_done_buf  = spc471_inst_done;
wire [63:0]                      pc_w471_buf           = pc_w471;


wire                             spc472_inst_done_buf  = spc472_inst_done;
wire [63:0]                      pc_w472_buf           = pc_w472;


wire                             spc473_inst_done_buf  = spc473_inst_done;
wire [63:0]                      pc_w473_buf           = pc_w473;


wire                             spc474_inst_done_buf  = spc474_inst_done;
wire [63:0]                      pc_w474_buf           = pc_w474;


wire                             spc475_inst_done_buf  = spc475_inst_done;
wire [63:0]                      pc_w475_buf           = pc_w475;


wire                             spc476_inst_done_buf  = spc476_inst_done;
wire [63:0]                      pc_w476_buf           = pc_w476;


wire                             spc477_inst_done_buf  = spc477_inst_done;
wire [63:0]                      pc_w477_buf           = pc_w477;


wire                             spc478_inst_done_buf  = spc478_inst_done;
wire [63:0]                      pc_w478_buf           = pc_w478;


wire                             spc479_inst_done_buf  = spc479_inst_done;
wire [63:0]                      pc_w479_buf           = pc_w479;


wire                             spc480_inst_done_buf  = spc480_inst_done;
wire [63:0]                      pc_w480_buf           = pc_w480;


wire                             spc481_inst_done_buf  = spc481_inst_done;
wire [63:0]                      pc_w481_buf           = pc_w481;


wire                             spc482_inst_done_buf  = spc482_inst_done;
wire [63:0]                      pc_w482_buf           = pc_w482;


wire                             spc483_inst_done_buf  = spc483_inst_done;
wire [63:0]                      pc_w483_buf           = pc_w483;


wire                             spc484_inst_done_buf  = spc484_inst_done;
wire [63:0]                      pc_w484_buf           = pc_w484;


wire                             spc485_inst_done_buf  = spc485_inst_done;
wire [63:0]                      pc_w485_buf           = pc_w485;


wire                             spc486_inst_done_buf  = spc486_inst_done;
wire [63:0]                      pc_w486_buf           = pc_w486;


wire                             spc487_inst_done_buf  = spc487_inst_done;
wire [63:0]                      pc_w487_buf           = pc_w487;


wire                             spc488_inst_done_buf  = spc488_inst_done;
wire [63:0]                      pc_w488_buf           = pc_w488;


wire                             spc489_inst_done_buf  = spc489_inst_done;
wire [63:0]                      pc_w489_buf           = pc_w489;


wire                             spc490_inst_done_buf  = spc490_inst_done;
wire [63:0]                      pc_w490_buf           = pc_w490;


wire                             spc491_inst_done_buf  = spc491_inst_done;
wire [63:0]                      pc_w491_buf           = pc_w491;


wire                             spc492_inst_done_buf  = spc492_inst_done;
wire [63:0]                      pc_w492_buf           = pc_w492;


wire                             spc493_inst_done_buf  = spc493_inst_done;
wire [63:0]                      pc_w493_buf           = pc_w493;


wire                             spc494_inst_done_buf  = spc494_inst_done;
wire [63:0]                      pc_w494_buf           = pc_w494;


wire                             spc495_inst_done_buf  = spc495_inst_done;
wire [63:0]                      pc_w495_buf           = pc_w495;


wire                             spc496_inst_done_buf  = spc496_inst_done;
wire [63:0]                      pc_w496_buf           = pc_w496;


wire                             spc497_inst_done_buf  = spc497_inst_done;
wire [63:0]                      pc_w497_buf           = pc_w497;


wire                             spc498_inst_done_buf  = spc498_inst_done;
wire [63:0]                      pc_w498_buf           = pc_w498;


wire                             spc499_inst_done_buf  = spc499_inst_done;
wire [63:0]                      pc_w499_buf           = pc_w499;


wire                             spc500_inst_done_buf  = spc500_inst_done;
wire [63:0]                      pc_w500_buf           = pc_w500;


wire                             spc501_inst_done_buf  = spc501_inst_done;
wire [63:0]                      pc_w501_buf           = pc_w501;


wire                             spc502_inst_done_buf  = spc502_inst_done;
wire [63:0]                      pc_w502_buf           = pc_w502;


wire                             spc503_inst_done_buf  = spc503_inst_done;
wire [63:0]                      pc_w503_buf           = pc_w503;


wire                             spc504_inst_done_buf  = spc504_inst_done;
wire [63:0]                      pc_w504_buf           = pc_w504;


wire                             spc505_inst_done_buf  = spc505_inst_done;
wire [63:0]                      pc_w505_buf           = pc_w505;


wire                             spc506_inst_done_buf  = spc506_inst_done;
wire [63:0]                      pc_w506_buf           = pc_w506;


wire                             spc507_inst_done_buf  = spc507_inst_done;
wire [63:0]                      pc_w507_buf           = pc_w507;


wire                             spc508_inst_done_buf  = spc508_inst_done;
wire [63:0]                      pc_w508_buf           = pc_w508;


wire                             spc509_inst_done_buf  = spc509_inst_done;
wire [63:0]                      pc_w509_buf           = pc_w509;


wire                             spc510_inst_done_buf  = spc510_inst_done;
wire [63:0]                      pc_w510_buf           = pc_w510;


wire                             spc511_inst_done_buf  = spc511_inst_done;
wire [63:0]                      pc_w511_buf           = pc_w511;


wire                             spc512_inst_done_buf  = spc512_inst_done;
wire [63:0]                      pc_w512_buf           = pc_w512;


wire                             spc513_inst_done_buf  = spc513_inst_done;
wire [63:0]                      pc_w513_buf           = pc_w513;


wire                             spc514_inst_done_buf  = spc514_inst_done;
wire [63:0]                      pc_w514_buf           = pc_w514;


wire                             spc515_inst_done_buf  = spc515_inst_done;
wire [63:0]                      pc_w515_buf           = pc_w515;


wire                             spc516_inst_done_buf  = spc516_inst_done;
wire [63:0]                      pc_w516_buf           = pc_w516;


wire                             spc517_inst_done_buf  = spc517_inst_done;
wire [63:0]                      pc_w517_buf           = pc_w517;


wire                             spc518_inst_done_buf  = spc518_inst_done;
wire [63:0]                      pc_w518_buf           = pc_w518;


wire                             spc519_inst_done_buf  = spc519_inst_done;
wire [63:0]                      pc_w519_buf           = pc_w519;


wire                             spc520_inst_done_buf  = spc520_inst_done;
wire [63:0]                      pc_w520_buf           = pc_w520;


wire                             spc521_inst_done_buf  = spc521_inst_done;
wire [63:0]                      pc_w521_buf           = pc_w521;


wire                             spc522_inst_done_buf  = spc522_inst_done;
wire [63:0]                      pc_w522_buf           = pc_w522;


wire                             spc523_inst_done_buf  = spc523_inst_done;
wire [63:0]                      pc_w523_buf           = pc_w523;


wire                             spc524_inst_done_buf  = spc524_inst_done;
wire [63:0]                      pc_w524_buf           = pc_w524;


wire                             spc525_inst_done_buf  = spc525_inst_done;
wire [63:0]                      pc_w525_buf           = pc_w525;


wire                             spc526_inst_done_buf  = spc526_inst_done;
wire [63:0]                      pc_w526_buf           = pc_w526;


wire                             spc527_inst_done_buf  = spc527_inst_done;
wire [63:0]                      pc_w527_buf           = pc_w527;


wire                             spc528_inst_done_buf  = spc528_inst_done;
wire [63:0]                      pc_w528_buf           = pc_w528;


wire                             spc529_inst_done_buf  = spc529_inst_done;
wire [63:0]                      pc_w529_buf           = pc_w529;


wire                             spc530_inst_done_buf  = spc530_inst_done;
wire [63:0]                      pc_w530_buf           = pc_w530;


wire                             spc531_inst_done_buf  = spc531_inst_done;
wire [63:0]                      pc_w531_buf           = pc_w531;


wire                             spc532_inst_done_buf  = spc532_inst_done;
wire [63:0]                      pc_w532_buf           = pc_w532;


wire                             spc533_inst_done_buf  = spc533_inst_done;
wire [63:0]                      pc_w533_buf           = pc_w533;


wire                             spc534_inst_done_buf  = spc534_inst_done;
wire [63:0]                      pc_w534_buf           = pc_w534;


wire                             spc535_inst_done_buf  = spc535_inst_done;
wire [63:0]                      pc_w535_buf           = pc_w535;


wire                             spc536_inst_done_buf  = spc536_inst_done;
wire [63:0]                      pc_w536_buf           = pc_w536;


wire                             spc537_inst_done_buf  = spc537_inst_done;
wire [63:0]                      pc_w537_buf           = pc_w537;


wire                             spc538_inst_done_buf  = spc538_inst_done;
wire [63:0]                      pc_w538_buf           = pc_w538;


wire                             spc539_inst_done_buf  = spc539_inst_done;
wire [63:0]                      pc_w539_buf           = pc_w539;


wire                             spc540_inst_done_buf  = spc540_inst_done;
wire [63:0]                      pc_w540_buf           = pc_w540;


wire                             spc541_inst_done_buf  = spc541_inst_done;
wire [63:0]                      pc_w541_buf           = pc_w541;


wire                             spc542_inst_done_buf  = spc542_inst_done;
wire [63:0]                      pc_w542_buf           = pc_w542;


wire                             spc543_inst_done_buf  = spc543_inst_done;
wire [63:0]                      pc_w543_buf           = pc_w543;


wire                             spc544_inst_done_buf  = spc544_inst_done;
wire [63:0]                      pc_w544_buf           = pc_w544;


wire                             spc545_inst_done_buf  = spc545_inst_done;
wire [63:0]                      pc_w545_buf           = pc_w545;


wire                             spc546_inst_done_buf  = spc546_inst_done;
wire [63:0]                      pc_w546_buf           = pc_w546;


wire                             spc547_inst_done_buf  = spc547_inst_done;
wire [63:0]                      pc_w547_buf           = pc_w547;


wire                             spc548_inst_done_buf  = spc548_inst_done;
wire [63:0]                      pc_w548_buf           = pc_w548;


wire                             spc549_inst_done_buf  = spc549_inst_done;
wire [63:0]                      pc_w549_buf           = pc_w549;


wire                             spc550_inst_done_buf  = spc550_inst_done;
wire [63:0]                      pc_w550_buf           = pc_w550;


wire                             spc551_inst_done_buf  = spc551_inst_done;
wire [63:0]                      pc_w551_buf           = pc_w551;


wire                             spc552_inst_done_buf  = spc552_inst_done;
wire [63:0]                      pc_w552_buf           = pc_w552;


wire                             spc553_inst_done_buf  = spc553_inst_done;
wire [63:0]                      pc_w553_buf           = pc_w553;


wire                             spc554_inst_done_buf  = spc554_inst_done;
wire [63:0]                      pc_w554_buf           = pc_w554;


wire                             spc555_inst_done_buf  = spc555_inst_done;
wire [63:0]                      pc_w555_buf           = pc_w555;


wire                             spc556_inst_done_buf  = spc556_inst_done;
wire [63:0]                      pc_w556_buf           = pc_w556;


wire                             spc557_inst_done_buf  = spc557_inst_done;
wire [63:0]                      pc_w557_buf           = pc_w557;


wire                             spc558_inst_done_buf  = spc558_inst_done;
wire [63:0]                      pc_w558_buf           = pc_w558;


wire                             spc559_inst_done_buf  = spc559_inst_done;
wire [63:0]                      pc_w559_buf           = pc_w559;


wire                             spc560_inst_done_buf  = spc560_inst_done;
wire [63:0]                      pc_w560_buf           = pc_w560;


wire                             spc561_inst_done_buf  = spc561_inst_done;
wire [63:0]                      pc_w561_buf           = pc_w561;


wire                             spc562_inst_done_buf  = spc562_inst_done;
wire [63:0]                      pc_w562_buf           = pc_w562;


wire                             spc563_inst_done_buf  = spc563_inst_done;
wire [63:0]                      pc_w563_buf           = pc_w563;


wire                             spc564_inst_done_buf  = spc564_inst_done;
wire [63:0]                      pc_w564_buf           = pc_w564;


wire                             spc565_inst_done_buf  = spc565_inst_done;
wire [63:0]                      pc_w565_buf           = pc_w565;


wire                             spc566_inst_done_buf  = spc566_inst_done;
wire [63:0]                      pc_w566_buf           = pc_w566;


wire                             spc567_inst_done_buf  = spc567_inst_done;
wire [63:0]                      pc_w567_buf           = pc_w567;


wire                             spc568_inst_done_buf  = spc568_inst_done;
wire [63:0]                      pc_w568_buf           = pc_w568;


wire                             spc569_inst_done_buf  = spc569_inst_done;
wire [63:0]                      pc_w569_buf           = pc_w569;


wire                             spc570_inst_done_buf  = spc570_inst_done;
wire [63:0]                      pc_w570_buf           = pc_w570;


wire                             spc571_inst_done_buf  = spc571_inst_done;
wire [63:0]                      pc_w571_buf           = pc_w571;


wire                             spc572_inst_done_buf  = spc572_inst_done;
wire [63:0]                      pc_w572_buf           = pc_w572;


wire                             spc573_inst_done_buf  = spc573_inst_done;
wire [63:0]                      pc_w573_buf           = pc_w573;


wire                             spc574_inst_done_buf  = spc574_inst_done;
wire [63:0]                      pc_w574_buf           = pc_w574;


wire                             spc575_inst_done_buf  = spc575_inst_done;
wire [63:0]                      pc_w575_buf           = pc_w575;


wire                             spc576_inst_done_buf  = spc576_inst_done;
wire [63:0]                      pc_w576_buf           = pc_w576;


wire                             spc577_inst_done_buf  = spc577_inst_done;
wire [63:0]                      pc_w577_buf           = pc_w577;


wire                             spc578_inst_done_buf  = spc578_inst_done;
wire [63:0]                      pc_w578_buf           = pc_w578;


wire                             spc579_inst_done_buf  = spc579_inst_done;
wire [63:0]                      pc_w579_buf           = pc_w579;


wire                             spc580_inst_done_buf  = spc580_inst_done;
wire [63:0]                      pc_w580_buf           = pc_w580;


wire                             spc581_inst_done_buf  = spc581_inst_done;
wire [63:0]                      pc_w581_buf           = pc_w581;


wire                             spc582_inst_done_buf  = spc582_inst_done;
wire [63:0]                      pc_w582_buf           = pc_w582;


wire                             spc583_inst_done_buf  = spc583_inst_done;
wire [63:0]                      pc_w583_buf           = pc_w583;


wire                             spc584_inst_done_buf  = spc584_inst_done;
wire [63:0]                      pc_w584_buf           = pc_w584;


wire                             spc585_inst_done_buf  = spc585_inst_done;
wire [63:0]                      pc_w585_buf           = pc_w585;


wire                             spc586_inst_done_buf  = spc586_inst_done;
wire [63:0]                      pc_w586_buf           = pc_w586;


wire                             spc587_inst_done_buf  = spc587_inst_done;
wire [63:0]                      pc_w587_buf           = pc_w587;


wire                             spc588_inst_done_buf  = spc588_inst_done;
wire [63:0]                      pc_w588_buf           = pc_w588;


wire                             spc589_inst_done_buf  = spc589_inst_done;
wire [63:0]                      pc_w589_buf           = pc_w589;


wire                             spc590_inst_done_buf  = spc590_inst_done;
wire [63:0]                      pc_w590_buf           = pc_w590;


wire                             spc591_inst_done_buf  = spc591_inst_done;
wire [63:0]                      pc_w591_buf           = pc_w591;


wire                             spc592_inst_done_buf  = spc592_inst_done;
wire [63:0]                      pc_w592_buf           = pc_w592;


wire                             spc593_inst_done_buf  = spc593_inst_done;
wire [63:0]                      pc_w593_buf           = pc_w593;


wire                             spc594_inst_done_buf  = spc594_inst_done;
wire [63:0]                      pc_w594_buf           = pc_w594;


wire                             spc595_inst_done_buf  = spc595_inst_done;
wire [63:0]                      pc_w595_buf           = pc_w595;


wire                             spc596_inst_done_buf  = spc596_inst_done;
wire [63:0]                      pc_w596_buf           = pc_w596;


wire                             spc597_inst_done_buf  = spc597_inst_done;
wire [63:0]                      pc_w597_buf           = pc_w597;


wire                             spc598_inst_done_buf  = spc598_inst_done;
wire [63:0]                      pc_w598_buf           = pc_w598;


wire                             spc599_inst_done_buf  = spc599_inst_done;
wire [63:0]                      pc_w599_buf           = pc_w599;


wire                             spc600_inst_done_buf  = spc600_inst_done;
wire [63:0]                      pc_w600_buf           = pc_w600;


wire                             spc601_inst_done_buf  = spc601_inst_done;
wire [63:0]                      pc_w601_buf           = pc_w601;


wire                             spc602_inst_done_buf  = spc602_inst_done;
wire [63:0]                      pc_w602_buf           = pc_w602;


wire                             spc603_inst_done_buf  = spc603_inst_done;
wire [63:0]                      pc_w603_buf           = pc_w603;


wire                             spc604_inst_done_buf  = spc604_inst_done;
wire [63:0]                      pc_w604_buf           = pc_w604;


wire                             spc605_inst_done_buf  = spc605_inst_done;
wire [63:0]                      pc_w605_buf           = pc_w605;


wire                             spc606_inst_done_buf  = spc606_inst_done;
wire [63:0]                      pc_w606_buf           = pc_w606;


wire                             spc607_inst_done_buf  = spc607_inst_done;
wire [63:0]                      pc_w607_buf           = pc_w607;


wire                             spc608_inst_done_buf  = spc608_inst_done;
wire [63:0]                      pc_w608_buf           = pc_w608;


wire                             spc609_inst_done_buf  = spc609_inst_done;
wire [63:0]                      pc_w609_buf           = pc_w609;


wire                             spc610_inst_done_buf  = spc610_inst_done;
wire [63:0]                      pc_w610_buf           = pc_w610;


wire                             spc611_inst_done_buf  = spc611_inst_done;
wire [63:0]                      pc_w611_buf           = pc_w611;


wire                             spc612_inst_done_buf  = spc612_inst_done;
wire [63:0]                      pc_w612_buf           = pc_w612;


wire                             spc613_inst_done_buf  = spc613_inst_done;
wire [63:0]                      pc_w613_buf           = pc_w613;


wire                             spc614_inst_done_buf  = spc614_inst_done;
wire [63:0]                      pc_w614_buf           = pc_w614;


wire                             spc615_inst_done_buf  = spc615_inst_done;
wire [63:0]                      pc_w615_buf           = pc_w615;


wire                             spc616_inst_done_buf  = spc616_inst_done;
wire [63:0]                      pc_w616_buf           = pc_w616;


wire                             spc617_inst_done_buf  = spc617_inst_done;
wire [63:0]                      pc_w617_buf           = pc_w617;


wire                             spc618_inst_done_buf  = spc618_inst_done;
wire [63:0]                      pc_w618_buf           = pc_w618;


wire                             spc619_inst_done_buf  = spc619_inst_done;
wire [63:0]                      pc_w619_buf           = pc_w619;


wire                             spc620_inst_done_buf  = spc620_inst_done;
wire [63:0]                      pc_w620_buf           = pc_w620;


wire                             spc621_inst_done_buf  = spc621_inst_done;
wire [63:0]                      pc_w621_buf           = pc_w621;


wire                             spc622_inst_done_buf  = spc622_inst_done;
wire [63:0]                      pc_w622_buf           = pc_w622;


wire                             spc623_inst_done_buf  = spc623_inst_done;
wire [63:0]                      pc_w623_buf           = pc_w623;


wire                             spc624_inst_done_buf  = spc624_inst_done;
wire [63:0]                      pc_w624_buf           = pc_w624;


wire                             spc625_inst_done_buf  = spc625_inst_done;
wire [63:0]                      pc_w625_buf           = pc_w625;


wire                             spc626_inst_done_buf  = spc626_inst_done;
wire [63:0]                      pc_w626_buf           = pc_w626;


wire                             spc627_inst_done_buf  = spc627_inst_done;
wire [63:0]                      pc_w627_buf           = pc_w627;


wire                             spc628_inst_done_buf  = spc628_inst_done;
wire [63:0]                      pc_w628_buf           = pc_w628;


wire                             spc629_inst_done_buf  = spc629_inst_done;
wire [63:0]                      pc_w629_buf           = pc_w629;


wire                             spc630_inst_done_buf  = spc630_inst_done;
wire [63:0]                      pc_w630_buf           = pc_w630;


wire                             spc631_inst_done_buf  = spc631_inst_done;
wire [63:0]                      pc_w631_buf           = pc_w631;


wire                             spc632_inst_done_buf  = spc632_inst_done;
wire [63:0]                      pc_w632_buf           = pc_w632;


wire                             spc633_inst_done_buf  = spc633_inst_done;
wire [63:0]                      pc_w633_buf           = pc_w633;


wire                             spc634_inst_done_buf  = spc634_inst_done;
wire [63:0]                      pc_w634_buf           = pc_w634;


wire                             spc635_inst_done_buf  = spc635_inst_done;
wire [63:0]                      pc_w635_buf           = pc_w635;


wire                             spc636_inst_done_buf  = spc636_inst_done;
wire [63:0]                      pc_w636_buf           = pc_w636;


wire                             spc637_inst_done_buf  = spc637_inst_done;
wire [63:0]                      pc_w637_buf           = pc_w637;


wire                             spc638_inst_done_buf  = spc638_inst_done;
wire [63:0]                      pc_w638_buf           = pc_w638;


wire                             spc639_inst_done_buf  = spc639_inst_done;
wire [63:0]                      pc_w639_buf           = pc_w639;


wire                             spc640_inst_done_buf  = spc640_inst_done;
wire [63:0]                      pc_w640_buf           = pc_w640;


wire                             spc641_inst_done_buf  = spc641_inst_done;
wire [63:0]                      pc_w641_buf           = pc_w641;


wire                             spc642_inst_done_buf  = spc642_inst_done;
wire [63:0]                      pc_w642_buf           = pc_w642;


wire                             spc643_inst_done_buf  = spc643_inst_done;
wire [63:0]                      pc_w643_buf           = pc_w643;


wire                             spc644_inst_done_buf  = spc644_inst_done;
wire [63:0]                      pc_w644_buf           = pc_w644;


wire                             spc645_inst_done_buf  = spc645_inst_done;
wire [63:0]                      pc_w645_buf           = pc_w645;


wire                             spc646_inst_done_buf  = spc646_inst_done;
wire [63:0]                      pc_w646_buf           = pc_w646;


wire                             spc647_inst_done_buf  = spc647_inst_done;
wire [63:0]                      pc_w647_buf           = pc_w647;


wire                             spc648_inst_done_buf  = spc648_inst_done;
wire [63:0]                      pc_w648_buf           = pc_w648;


wire                             spc649_inst_done_buf  = spc649_inst_done;
wire [63:0]                      pc_w649_buf           = pc_w649;


wire                             spc650_inst_done_buf  = spc650_inst_done;
wire [63:0]                      pc_w650_buf           = pc_w650;


wire                             spc651_inst_done_buf  = spc651_inst_done;
wire [63:0]                      pc_w651_buf           = pc_w651;


wire                             spc652_inst_done_buf  = spc652_inst_done;
wire [63:0]                      pc_w652_buf           = pc_w652;


wire                             spc653_inst_done_buf  = spc653_inst_done;
wire [63:0]                      pc_w653_buf           = pc_w653;


wire                             spc654_inst_done_buf  = spc654_inst_done;
wire [63:0]                      pc_w654_buf           = pc_w654;


wire                             spc655_inst_done_buf  = spc655_inst_done;
wire [63:0]                      pc_w655_buf           = pc_w655;


wire                             spc656_inst_done_buf  = spc656_inst_done;
wire [63:0]                      pc_w656_buf           = pc_w656;


wire                             spc657_inst_done_buf  = spc657_inst_done;
wire [63:0]                      pc_w657_buf           = pc_w657;


wire                             spc658_inst_done_buf  = spc658_inst_done;
wire [63:0]                      pc_w658_buf           = pc_w658;


wire                             spc659_inst_done_buf  = spc659_inst_done;
wire [63:0]                      pc_w659_buf           = pc_w659;


wire                             spc660_inst_done_buf  = spc660_inst_done;
wire [63:0]                      pc_w660_buf           = pc_w660;


wire                             spc661_inst_done_buf  = spc661_inst_done;
wire [63:0]                      pc_w661_buf           = pc_w661;


wire                             spc662_inst_done_buf  = spc662_inst_done;
wire [63:0]                      pc_w662_buf           = pc_w662;


wire                             spc663_inst_done_buf  = spc663_inst_done;
wire [63:0]                      pc_w663_buf           = pc_w663;


wire                             spc664_inst_done_buf  = spc664_inst_done;
wire [63:0]                      pc_w664_buf           = pc_w664;


wire                             spc665_inst_done_buf  = spc665_inst_done;
wire [63:0]                      pc_w665_buf           = pc_w665;


wire                             spc666_inst_done_buf  = spc666_inst_done;
wire [63:0]                      pc_w666_buf           = pc_w666;


wire                             spc667_inst_done_buf  = spc667_inst_done;
wire [63:0]                      pc_w667_buf           = pc_w667;


wire                             spc668_inst_done_buf  = spc668_inst_done;
wire [63:0]                      pc_w668_buf           = pc_w668;


wire                             spc669_inst_done_buf  = spc669_inst_done;
wire [63:0]                      pc_w669_buf           = pc_w669;


wire                             spc670_inst_done_buf  = spc670_inst_done;
wire [63:0]                      pc_w670_buf           = pc_w670;


wire                             spc671_inst_done_buf  = spc671_inst_done;
wire [63:0]                      pc_w671_buf           = pc_w671;


wire                             spc672_inst_done_buf  = spc672_inst_done;
wire [63:0]                      pc_w672_buf           = pc_w672;


wire                             spc673_inst_done_buf  = spc673_inst_done;
wire [63:0]                      pc_w673_buf           = pc_w673;


wire                             spc674_inst_done_buf  = spc674_inst_done;
wire [63:0]                      pc_w674_buf           = pc_w674;


wire                             spc675_inst_done_buf  = spc675_inst_done;
wire [63:0]                      pc_w675_buf           = pc_w675;


wire                             spc676_inst_done_buf  = spc676_inst_done;
wire [63:0]                      pc_w676_buf           = pc_w676;


wire                             spc677_inst_done_buf  = spc677_inst_done;
wire [63:0]                      pc_w677_buf           = pc_w677;


wire                             spc678_inst_done_buf  = spc678_inst_done;
wire [63:0]                      pc_w678_buf           = pc_w678;


wire                             spc679_inst_done_buf  = spc679_inst_done;
wire [63:0]                      pc_w679_buf           = pc_w679;


wire                             spc680_inst_done_buf  = spc680_inst_done;
wire [63:0]                      pc_w680_buf           = pc_w680;


wire                             spc681_inst_done_buf  = spc681_inst_done;
wire [63:0]                      pc_w681_buf           = pc_w681;


wire                             spc682_inst_done_buf  = spc682_inst_done;
wire [63:0]                      pc_w682_buf           = pc_w682;


wire                             spc683_inst_done_buf  = spc683_inst_done;
wire [63:0]                      pc_w683_buf           = pc_w683;


wire                             spc684_inst_done_buf  = spc684_inst_done;
wire [63:0]                      pc_w684_buf           = pc_w684;


wire                             spc685_inst_done_buf  = spc685_inst_done;
wire [63:0]                      pc_w685_buf           = pc_w685;


wire                             spc686_inst_done_buf  = spc686_inst_done;
wire [63:0]                      pc_w686_buf           = pc_w686;


wire                             spc687_inst_done_buf  = spc687_inst_done;
wire [63:0]                      pc_w687_buf           = pc_w687;


wire                             spc688_inst_done_buf  = spc688_inst_done;
wire [63:0]                      pc_w688_buf           = pc_w688;


wire                             spc689_inst_done_buf  = spc689_inst_done;
wire [63:0]                      pc_w689_buf           = pc_w689;


wire                             spc690_inst_done_buf  = spc690_inst_done;
wire [63:0]                      pc_w690_buf           = pc_w690;


wire                             spc691_inst_done_buf  = spc691_inst_done;
wire [63:0]                      pc_w691_buf           = pc_w691;


wire                             spc692_inst_done_buf  = spc692_inst_done;
wire [63:0]                      pc_w692_buf           = pc_w692;


wire                             spc693_inst_done_buf  = spc693_inst_done;
wire [63:0]                      pc_w693_buf           = pc_w693;


wire                             spc694_inst_done_buf  = spc694_inst_done;
wire [63:0]                      pc_w694_buf           = pc_w694;


wire                             spc695_inst_done_buf  = spc695_inst_done;
wire [63:0]                      pc_w695_buf           = pc_w695;


wire                             spc696_inst_done_buf  = spc696_inst_done;
wire [63:0]                      pc_w696_buf           = pc_w696;


wire                             spc697_inst_done_buf  = spc697_inst_done;
wire [63:0]                      pc_w697_buf           = pc_w697;


wire                             spc698_inst_done_buf  = spc698_inst_done;
wire [63:0]                      pc_w698_buf           = pc_w698;


wire                             spc699_inst_done_buf  = spc699_inst_done;
wire [63:0]                      pc_w699_buf           = pc_w699;


wire                             spc700_inst_done_buf  = spc700_inst_done;
wire [63:0]                      pc_w700_buf           = pc_w700;


wire                             spc701_inst_done_buf  = spc701_inst_done;
wire [63:0]                      pc_w701_buf           = pc_w701;


wire                             spc702_inst_done_buf  = spc702_inst_done;
wire [63:0]                      pc_w702_buf           = pc_w702;


wire                             spc703_inst_done_buf  = spc703_inst_done;
wire [63:0]                      pc_w703_buf           = pc_w703;


wire                             spc704_inst_done_buf  = spc704_inst_done;
wire [63:0]                      pc_w704_buf           = pc_w704;


wire                             spc705_inst_done_buf  = spc705_inst_done;
wire [63:0]                      pc_w705_buf           = pc_w705;


wire                             spc706_inst_done_buf  = spc706_inst_done;
wire [63:0]                      pc_w706_buf           = pc_w706;


wire                             spc707_inst_done_buf  = spc707_inst_done;
wire [63:0]                      pc_w707_buf           = pc_w707;


wire                             spc708_inst_done_buf  = spc708_inst_done;
wire [63:0]                      pc_w708_buf           = pc_w708;


wire                             spc709_inst_done_buf  = spc709_inst_done;
wire [63:0]                      pc_w709_buf           = pc_w709;


wire                             spc710_inst_done_buf  = spc710_inst_done;
wire [63:0]                      pc_w710_buf           = pc_w710;


wire                             spc711_inst_done_buf  = spc711_inst_done;
wire [63:0]                      pc_w711_buf           = pc_w711;


wire                             spc712_inst_done_buf  = spc712_inst_done;
wire [63:0]                      pc_w712_buf           = pc_w712;


wire                             spc713_inst_done_buf  = spc713_inst_done;
wire [63:0]                      pc_w713_buf           = pc_w713;


wire                             spc714_inst_done_buf  = spc714_inst_done;
wire [63:0]                      pc_w714_buf           = pc_w714;


wire                             spc715_inst_done_buf  = spc715_inst_done;
wire [63:0]                      pc_w715_buf           = pc_w715;


wire                             spc716_inst_done_buf  = spc716_inst_done;
wire [63:0]                      pc_w716_buf           = pc_w716;


wire                             spc717_inst_done_buf  = spc717_inst_done;
wire [63:0]                      pc_w717_buf           = pc_w717;


wire                             spc718_inst_done_buf  = spc718_inst_done;
wire [63:0]                      pc_w718_buf           = pc_w718;


wire                             spc719_inst_done_buf  = spc719_inst_done;
wire [63:0]                      pc_w719_buf           = pc_w719;


wire                             spc720_inst_done_buf  = spc720_inst_done;
wire [63:0]                      pc_w720_buf           = pc_w720;


wire                             spc721_inst_done_buf  = spc721_inst_done;
wire [63:0]                      pc_w721_buf           = pc_w721;


wire                             spc722_inst_done_buf  = spc722_inst_done;
wire [63:0]                      pc_w722_buf           = pc_w722;


wire                             spc723_inst_done_buf  = spc723_inst_done;
wire [63:0]                      pc_w723_buf           = pc_w723;


wire                             spc724_inst_done_buf  = spc724_inst_done;
wire [63:0]                      pc_w724_buf           = pc_w724;


wire                             spc725_inst_done_buf  = spc725_inst_done;
wire [63:0]                      pc_w725_buf           = pc_w725;


wire                             spc726_inst_done_buf  = spc726_inst_done;
wire [63:0]                      pc_w726_buf           = pc_w726;


wire                             spc727_inst_done_buf  = spc727_inst_done;
wire [63:0]                      pc_w727_buf           = pc_w727;


wire                             spc728_inst_done_buf  = spc728_inst_done;
wire [63:0]                      pc_w728_buf           = pc_w728;


wire                             spc729_inst_done_buf  = spc729_inst_done;
wire [63:0]                      pc_w729_buf           = pc_w729;


wire                             spc730_inst_done_buf  = spc730_inst_done;
wire [63:0]                      pc_w730_buf           = pc_w730;


wire                             spc731_inst_done_buf  = spc731_inst_done;
wire [63:0]                      pc_w731_buf           = pc_w731;


wire                             spc732_inst_done_buf  = spc732_inst_done;
wire [63:0]                      pc_w732_buf           = pc_w732;


wire                             spc733_inst_done_buf  = spc733_inst_done;
wire [63:0]                      pc_w733_buf           = pc_w733;


wire                             spc734_inst_done_buf  = spc734_inst_done;
wire [63:0]                      pc_w734_buf           = pc_w734;


wire                             spc735_inst_done_buf  = spc735_inst_done;
wire [63:0]                      pc_w735_buf           = pc_w735;


wire                             spc736_inst_done_buf  = spc736_inst_done;
wire [63:0]                      pc_w736_buf           = pc_w736;


wire                             spc737_inst_done_buf  = spc737_inst_done;
wire [63:0]                      pc_w737_buf           = pc_w737;


wire                             spc738_inst_done_buf  = spc738_inst_done;
wire [63:0]                      pc_w738_buf           = pc_w738;


wire                             spc739_inst_done_buf  = spc739_inst_done;
wire [63:0]                      pc_w739_buf           = pc_w739;


wire                             spc740_inst_done_buf  = spc740_inst_done;
wire [63:0]                      pc_w740_buf           = pc_w740;


wire                             spc741_inst_done_buf  = spc741_inst_done;
wire [63:0]                      pc_w741_buf           = pc_w741;


wire                             spc742_inst_done_buf  = spc742_inst_done;
wire [63:0]                      pc_w742_buf           = pc_w742;


wire                             spc743_inst_done_buf  = spc743_inst_done;
wire [63:0]                      pc_w743_buf           = pc_w743;


wire                             spc744_inst_done_buf  = spc744_inst_done;
wire [63:0]                      pc_w744_buf           = pc_w744;


wire                             spc745_inst_done_buf  = spc745_inst_done;
wire [63:0]                      pc_w745_buf           = pc_w745;


wire                             spc746_inst_done_buf  = spc746_inst_done;
wire [63:0]                      pc_w746_buf           = pc_w746;


wire                             spc747_inst_done_buf  = spc747_inst_done;
wire [63:0]                      pc_w747_buf           = pc_w747;


wire                             spc748_inst_done_buf  = spc748_inst_done;
wire [63:0]                      pc_w748_buf           = pc_w748;


wire                             spc749_inst_done_buf  = spc749_inst_done;
wire [63:0]                      pc_w749_buf           = pc_w749;


wire                             spc750_inst_done_buf  = spc750_inst_done;
wire [63:0]                      pc_w750_buf           = pc_w750;


wire                             spc751_inst_done_buf  = spc751_inst_done;
wire [63:0]                      pc_w751_buf           = pc_w751;


wire                             spc752_inst_done_buf  = spc752_inst_done;
wire [63:0]                      pc_w752_buf           = pc_w752;


wire                             spc753_inst_done_buf  = spc753_inst_done;
wire [63:0]                      pc_w753_buf           = pc_w753;


wire                             spc754_inst_done_buf  = spc754_inst_done;
wire [63:0]                      pc_w754_buf           = pc_w754;


wire                             spc755_inst_done_buf  = spc755_inst_done;
wire [63:0]                      pc_w755_buf           = pc_w755;


wire                             spc756_inst_done_buf  = spc756_inst_done;
wire [63:0]                      pc_w756_buf           = pc_w756;


wire                             spc757_inst_done_buf  = spc757_inst_done;
wire [63:0]                      pc_w757_buf           = pc_w757;


wire                             spc758_inst_done_buf  = spc758_inst_done;
wire [63:0]                      pc_w758_buf           = pc_w758;


wire                             spc759_inst_done_buf  = spc759_inst_done;
wire [63:0]                      pc_w759_buf           = pc_w759;


wire                             spc760_inst_done_buf  = spc760_inst_done;
wire [63:0]                      pc_w760_buf           = pc_w760;


wire                             spc761_inst_done_buf  = spc761_inst_done;
wire [63:0]                      pc_w761_buf           = pc_w761;


wire                             spc762_inst_done_buf  = spc762_inst_done;
wire [63:0]                      pc_w762_buf           = pc_w762;


wire                             spc763_inst_done_buf  = spc763_inst_done;
wire [63:0]                      pc_w763_buf           = pc_w763;


wire                             spc764_inst_done_buf  = spc764_inst_done;
wire [63:0]                      pc_w764_buf           = pc_w764;


wire                             spc765_inst_done_buf  = spc765_inst_done;
wire [63:0]                      pc_w765_buf           = pc_w765;


wire                             spc766_inst_done_buf  = spc766_inst_done;
wire [63:0]                      pc_w766_buf           = pc_w766;


wire                             spc767_inst_done_buf  = spc767_inst_done;
wire [63:0]                      pc_w767_buf           = pc_w767;


wire                             spc768_inst_done_buf  = spc768_inst_done;
wire [63:0]                      pc_w768_buf           = pc_w768;


wire                             spc769_inst_done_buf  = spc769_inst_done;
wire [63:0]                      pc_w769_buf           = pc_w769;


wire                             spc770_inst_done_buf  = spc770_inst_done;
wire [63:0]                      pc_w770_buf           = pc_w770;


wire                             spc771_inst_done_buf  = spc771_inst_done;
wire [63:0]                      pc_w771_buf           = pc_w771;


wire                             spc772_inst_done_buf  = spc772_inst_done;
wire [63:0]                      pc_w772_buf           = pc_w772;


wire                             spc773_inst_done_buf  = spc773_inst_done;
wire [63:0]                      pc_w773_buf           = pc_w773;


wire                             spc774_inst_done_buf  = spc774_inst_done;
wire [63:0]                      pc_w774_buf           = pc_w774;


wire                             spc775_inst_done_buf  = spc775_inst_done;
wire [63:0]                      pc_w775_buf           = pc_w775;


wire                             spc776_inst_done_buf  = spc776_inst_done;
wire [63:0]                      pc_w776_buf           = pc_w776;


wire                             spc777_inst_done_buf  = spc777_inst_done;
wire [63:0]                      pc_w777_buf           = pc_w777;


wire                             spc778_inst_done_buf  = spc778_inst_done;
wire [63:0]                      pc_w778_buf           = pc_w778;


wire                             spc779_inst_done_buf  = spc779_inst_done;
wire [63:0]                      pc_w779_buf           = pc_w779;


wire                             spc780_inst_done_buf  = spc780_inst_done;
wire [63:0]                      pc_w780_buf           = pc_w780;


wire                             spc781_inst_done_buf  = spc781_inst_done;
wire [63:0]                      pc_w781_buf           = pc_w781;


wire                             spc782_inst_done_buf  = spc782_inst_done;
wire [63:0]                      pc_w782_buf           = pc_w782;


wire                             spc783_inst_done_buf  = spc783_inst_done;
wire [63:0]                      pc_w783_buf           = pc_w783;


wire                             spc784_inst_done_buf  = spc784_inst_done;
wire [63:0]                      pc_w784_buf           = pc_w784;


wire                             spc785_inst_done_buf  = spc785_inst_done;
wire [63:0]                      pc_w785_buf           = pc_w785;


wire                             spc786_inst_done_buf  = spc786_inst_done;
wire [63:0]                      pc_w786_buf           = pc_w786;


wire                             spc787_inst_done_buf  = spc787_inst_done;
wire [63:0]                      pc_w787_buf           = pc_w787;


wire                             spc788_inst_done_buf  = spc788_inst_done;
wire [63:0]                      pc_w788_buf           = pc_w788;


wire                             spc789_inst_done_buf  = spc789_inst_done;
wire [63:0]                      pc_w789_buf           = pc_w789;


wire                             spc790_inst_done_buf  = spc790_inst_done;
wire [63:0]                      pc_w790_buf           = pc_w790;


wire                             spc791_inst_done_buf  = spc791_inst_done;
wire [63:0]                      pc_w791_buf           = pc_w791;


wire                             spc792_inst_done_buf  = spc792_inst_done;
wire [63:0]                      pc_w792_buf           = pc_w792;


wire                             spc793_inst_done_buf  = spc793_inst_done;
wire [63:0]                      pc_w793_buf           = pc_w793;


wire                             spc794_inst_done_buf  = spc794_inst_done;
wire [63:0]                      pc_w794_buf           = pc_w794;


wire                             spc795_inst_done_buf  = spc795_inst_done;
wire [63:0]                      pc_w795_buf           = pc_w795;


wire                             spc796_inst_done_buf  = spc796_inst_done;
wire [63:0]                      pc_w796_buf           = pc_w796;


wire                             spc797_inst_done_buf  = spc797_inst_done;
wire [63:0]                      pc_w797_buf           = pc_w797;


wire                             spc798_inst_done_buf  = spc798_inst_done;
wire [63:0]                      pc_w798_buf           = pc_w798;


wire                             spc799_inst_done_buf  = spc799_inst_done;
wire [63:0]                      pc_w799_buf           = pc_w799;


wire                             spc800_inst_done_buf  = spc800_inst_done;
wire [63:0]                      pc_w800_buf           = pc_w800;


wire                             spc801_inst_done_buf  = spc801_inst_done;
wire [63:0]                      pc_w801_buf           = pc_w801;


wire                             spc802_inst_done_buf  = spc802_inst_done;
wire [63:0]                      pc_w802_buf           = pc_w802;


wire                             spc803_inst_done_buf  = spc803_inst_done;
wire [63:0]                      pc_w803_buf           = pc_w803;


wire                             spc804_inst_done_buf  = spc804_inst_done;
wire [63:0]                      pc_w804_buf           = pc_w804;


wire                             spc805_inst_done_buf  = spc805_inst_done;
wire [63:0]                      pc_w805_buf           = pc_w805;


wire                             spc806_inst_done_buf  = spc806_inst_done;
wire [63:0]                      pc_w806_buf           = pc_w806;


wire                             spc807_inst_done_buf  = spc807_inst_done;
wire [63:0]                      pc_w807_buf           = pc_w807;


wire                             spc808_inst_done_buf  = spc808_inst_done;
wire [63:0]                      pc_w808_buf           = pc_w808;


wire                             spc809_inst_done_buf  = spc809_inst_done;
wire [63:0]                      pc_w809_buf           = pc_w809;


wire                             spc810_inst_done_buf  = spc810_inst_done;
wire [63:0]                      pc_w810_buf           = pc_w810;


wire                             spc811_inst_done_buf  = spc811_inst_done;
wire [63:0]                      pc_w811_buf           = pc_w811;


wire                             spc812_inst_done_buf  = spc812_inst_done;
wire [63:0]                      pc_w812_buf           = pc_w812;


wire                             spc813_inst_done_buf  = spc813_inst_done;
wire [63:0]                      pc_w813_buf           = pc_w813;


wire                             spc814_inst_done_buf  = spc814_inst_done;
wire [63:0]                      pc_w814_buf           = pc_w814;


wire                             spc815_inst_done_buf  = spc815_inst_done;
wire [63:0]                      pc_w815_buf           = pc_w815;


wire                             spc816_inst_done_buf  = spc816_inst_done;
wire [63:0]                      pc_w816_buf           = pc_w816;


wire                             spc817_inst_done_buf  = spc817_inst_done;
wire [63:0]                      pc_w817_buf           = pc_w817;


wire                             spc818_inst_done_buf  = spc818_inst_done;
wire [63:0]                      pc_w818_buf           = pc_w818;


wire                             spc819_inst_done_buf  = spc819_inst_done;
wire [63:0]                      pc_w819_buf           = pc_w819;


wire                             spc820_inst_done_buf  = spc820_inst_done;
wire [63:0]                      pc_w820_buf           = pc_w820;


wire                             spc821_inst_done_buf  = spc821_inst_done;
wire [63:0]                      pc_w821_buf           = pc_w821;


wire                             spc822_inst_done_buf  = spc822_inst_done;
wire [63:0]                      pc_w822_buf           = pc_w822;


wire                             spc823_inst_done_buf  = spc823_inst_done;
wire [63:0]                      pc_w823_buf           = pc_w823;


wire                             spc824_inst_done_buf  = spc824_inst_done;
wire [63:0]                      pc_w824_buf           = pc_w824;


wire                             spc825_inst_done_buf  = spc825_inst_done;
wire [63:0]                      pc_w825_buf           = pc_w825;


wire                             spc826_inst_done_buf  = spc826_inst_done;
wire [63:0]                      pc_w826_buf           = pc_w826;


wire                             spc827_inst_done_buf  = spc827_inst_done;
wire [63:0]                      pc_w827_buf           = pc_w827;


wire                             spc828_inst_done_buf  = spc828_inst_done;
wire [63:0]                      pc_w828_buf           = pc_w828;


wire                             spc829_inst_done_buf  = spc829_inst_done;
wire [63:0]                      pc_w829_buf           = pc_w829;


wire                             spc830_inst_done_buf  = spc830_inst_done;
wire [63:0]                      pc_w830_buf           = pc_w830;


wire                             spc831_inst_done_buf  = spc831_inst_done;
wire [63:0]                      pc_w831_buf           = pc_w831;


wire                             spc832_inst_done_buf  = spc832_inst_done;
wire [63:0]                      pc_w832_buf           = pc_w832;


wire                             spc833_inst_done_buf  = spc833_inst_done;
wire [63:0]                      pc_w833_buf           = pc_w833;


wire                             spc834_inst_done_buf  = spc834_inst_done;
wire [63:0]                      pc_w834_buf           = pc_w834;


wire                             spc835_inst_done_buf  = spc835_inst_done;
wire [63:0]                      pc_w835_buf           = pc_w835;


wire                             spc836_inst_done_buf  = spc836_inst_done;
wire [63:0]                      pc_w836_buf           = pc_w836;


wire                             spc837_inst_done_buf  = spc837_inst_done;
wire [63:0]                      pc_w837_buf           = pc_w837;


wire                             spc838_inst_done_buf  = spc838_inst_done;
wire [63:0]                      pc_w838_buf           = pc_w838;


wire                             spc839_inst_done_buf  = spc839_inst_done;
wire [63:0]                      pc_w839_buf           = pc_w839;


wire                             spc840_inst_done_buf  = spc840_inst_done;
wire [63:0]                      pc_w840_buf           = pc_w840;


wire                             spc841_inst_done_buf  = spc841_inst_done;
wire [63:0]                      pc_w841_buf           = pc_w841;


wire                             spc842_inst_done_buf  = spc842_inst_done;
wire [63:0]                      pc_w842_buf           = pc_w842;


wire                             spc843_inst_done_buf  = spc843_inst_done;
wire [63:0]                      pc_w843_buf           = pc_w843;


wire                             spc844_inst_done_buf  = spc844_inst_done;
wire [63:0]                      pc_w844_buf           = pc_w844;


wire                             spc845_inst_done_buf  = spc845_inst_done;
wire [63:0]                      pc_w845_buf           = pc_w845;


wire                             spc846_inst_done_buf  = spc846_inst_done;
wire [63:0]                      pc_w846_buf           = pc_w846;


wire                             spc847_inst_done_buf  = spc847_inst_done;
wire [63:0]                      pc_w847_buf           = pc_w847;


wire                             spc848_inst_done_buf  = spc848_inst_done;
wire [63:0]                      pc_w848_buf           = pc_w848;


wire                             spc849_inst_done_buf  = spc849_inst_done;
wire [63:0]                      pc_w849_buf           = pc_w849;


wire                             spc850_inst_done_buf  = spc850_inst_done;
wire [63:0]                      pc_w850_buf           = pc_w850;


wire                             spc851_inst_done_buf  = spc851_inst_done;
wire [63:0]                      pc_w851_buf           = pc_w851;


wire                             spc852_inst_done_buf  = spc852_inst_done;
wire [63:0]                      pc_w852_buf           = pc_w852;


wire                             spc853_inst_done_buf  = spc853_inst_done;
wire [63:0]                      pc_w853_buf           = pc_w853;


wire                             spc854_inst_done_buf  = spc854_inst_done;
wire [63:0]                      pc_w854_buf           = pc_w854;


wire                             spc855_inst_done_buf  = spc855_inst_done;
wire [63:0]                      pc_w855_buf           = pc_w855;


wire                             spc856_inst_done_buf  = spc856_inst_done;
wire [63:0]                      pc_w856_buf           = pc_w856;


wire                             spc857_inst_done_buf  = spc857_inst_done;
wire [63:0]                      pc_w857_buf           = pc_w857;


wire                             spc858_inst_done_buf  = spc858_inst_done;
wire [63:0]                      pc_w858_buf           = pc_w858;


wire                             spc859_inst_done_buf  = spc859_inst_done;
wire [63:0]                      pc_w859_buf           = pc_w859;


wire                             spc860_inst_done_buf  = spc860_inst_done;
wire [63:0]                      pc_w860_buf           = pc_w860;


wire                             spc861_inst_done_buf  = spc861_inst_done;
wire [63:0]                      pc_w861_buf           = pc_w861;


wire                             spc862_inst_done_buf  = spc862_inst_done;
wire [63:0]                      pc_w862_buf           = pc_w862;


wire                             spc863_inst_done_buf  = spc863_inst_done;
wire [63:0]                      pc_w863_buf           = pc_w863;


wire                             spc864_inst_done_buf  = spc864_inst_done;
wire [63:0]                      pc_w864_buf           = pc_w864;


wire                             spc865_inst_done_buf  = spc865_inst_done;
wire [63:0]                      pc_w865_buf           = pc_w865;


wire                             spc866_inst_done_buf  = spc866_inst_done;
wire [63:0]                      pc_w866_buf           = pc_w866;


wire                             spc867_inst_done_buf  = spc867_inst_done;
wire [63:0]                      pc_w867_buf           = pc_w867;


wire                             spc868_inst_done_buf  = spc868_inst_done;
wire [63:0]                      pc_w868_buf           = pc_w868;


wire                             spc869_inst_done_buf  = spc869_inst_done;
wire [63:0]                      pc_w869_buf           = pc_w869;


wire                             spc870_inst_done_buf  = spc870_inst_done;
wire [63:0]                      pc_w870_buf           = pc_w870;


wire                             spc871_inst_done_buf  = spc871_inst_done;
wire [63:0]                      pc_w871_buf           = pc_w871;


wire                             spc872_inst_done_buf  = spc872_inst_done;
wire [63:0]                      pc_w872_buf           = pc_w872;


wire                             spc873_inst_done_buf  = spc873_inst_done;
wire [63:0]                      pc_w873_buf           = pc_w873;


wire                             spc874_inst_done_buf  = spc874_inst_done;
wire [63:0]                      pc_w874_buf           = pc_w874;


wire                             spc875_inst_done_buf  = spc875_inst_done;
wire [63:0]                      pc_w875_buf           = pc_w875;


wire                             spc876_inst_done_buf  = spc876_inst_done;
wire [63:0]                      pc_w876_buf           = pc_w876;


wire                             spc877_inst_done_buf  = spc877_inst_done;
wire [63:0]                      pc_w877_buf           = pc_w877;


wire                             spc878_inst_done_buf  = spc878_inst_done;
wire [63:0]                      pc_w878_buf           = pc_w878;


wire                             spc879_inst_done_buf  = spc879_inst_done;
wire [63:0]                      pc_w879_buf           = pc_w879;


wire                             spc880_inst_done_buf  = spc880_inst_done;
wire [63:0]                      pc_w880_buf           = pc_w880;


wire                             spc881_inst_done_buf  = spc881_inst_done;
wire [63:0]                      pc_w881_buf           = pc_w881;


wire                             spc882_inst_done_buf  = spc882_inst_done;
wire [63:0]                      pc_w882_buf           = pc_w882;


wire                             spc883_inst_done_buf  = spc883_inst_done;
wire [63:0]                      pc_w883_buf           = pc_w883;


wire                             spc884_inst_done_buf  = spc884_inst_done;
wire [63:0]                      pc_w884_buf           = pc_w884;


wire                             spc885_inst_done_buf  = spc885_inst_done;
wire [63:0]                      pc_w885_buf           = pc_w885;


wire                             spc886_inst_done_buf  = spc886_inst_done;
wire [63:0]                      pc_w886_buf           = pc_w886;


wire                             spc887_inst_done_buf  = spc887_inst_done;
wire [63:0]                      pc_w887_buf           = pc_w887;


wire                             spc888_inst_done_buf  = spc888_inst_done;
wire [63:0]                      pc_w888_buf           = pc_w888;


wire                             spc889_inst_done_buf  = spc889_inst_done;
wire [63:0]                      pc_w889_buf           = pc_w889;


wire                             spc890_inst_done_buf  = spc890_inst_done;
wire [63:0]                      pc_w890_buf           = pc_w890;


wire                             spc891_inst_done_buf  = spc891_inst_done;
wire [63:0]                      pc_w891_buf           = pc_w891;


wire                             spc892_inst_done_buf  = spc892_inst_done;
wire [63:0]                      pc_w892_buf           = pc_w892;


wire                             spc893_inst_done_buf  = spc893_inst_done;
wire [63:0]                      pc_w893_buf           = pc_w893;


wire                             spc894_inst_done_buf  = spc894_inst_done;
wire [63:0]                      pc_w894_buf           = pc_w894;


wire                             spc895_inst_done_buf  = spc895_inst_done;
wire [63:0]                      pc_w895_buf           = pc_w895;


wire                             spc896_inst_done_buf  = spc896_inst_done;
wire [63:0]                      pc_w896_buf           = pc_w896;


wire                             spc897_inst_done_buf  = spc897_inst_done;
wire [63:0]                      pc_w897_buf           = pc_w897;


wire                             spc898_inst_done_buf  = spc898_inst_done;
wire [63:0]                      pc_w898_buf           = pc_w898;


wire                             spc899_inst_done_buf  = spc899_inst_done;
wire [63:0]                      pc_w899_buf           = pc_w899;


wire                             spc900_inst_done_buf  = spc900_inst_done;
wire [63:0]                      pc_w900_buf           = pc_w900;


wire                             spc901_inst_done_buf  = spc901_inst_done;
wire [63:0]                      pc_w901_buf           = pc_w901;


wire                             spc902_inst_done_buf  = spc902_inst_done;
wire [63:0]                      pc_w902_buf           = pc_w902;


wire                             spc903_inst_done_buf  = spc903_inst_done;
wire [63:0]                      pc_w903_buf           = pc_w903;


wire                             spc904_inst_done_buf  = spc904_inst_done;
wire [63:0]                      pc_w904_buf           = pc_w904;


wire                             spc905_inst_done_buf  = spc905_inst_done;
wire [63:0]                      pc_w905_buf           = pc_w905;


wire                             spc906_inst_done_buf  = spc906_inst_done;
wire [63:0]                      pc_w906_buf           = pc_w906;


wire                             spc907_inst_done_buf  = spc907_inst_done;
wire [63:0]                      pc_w907_buf           = pc_w907;


wire                             spc908_inst_done_buf  = spc908_inst_done;
wire [63:0]                      pc_w908_buf           = pc_w908;


wire                             spc909_inst_done_buf  = spc909_inst_done;
wire [63:0]                      pc_w909_buf           = pc_w909;


wire                             spc910_inst_done_buf  = spc910_inst_done;
wire [63:0]                      pc_w910_buf           = pc_w910;


wire                             spc911_inst_done_buf  = spc911_inst_done;
wire [63:0]                      pc_w911_buf           = pc_w911;


wire                             spc912_inst_done_buf  = spc912_inst_done;
wire [63:0]                      pc_w912_buf           = pc_w912;


wire                             spc913_inst_done_buf  = spc913_inst_done;
wire [63:0]                      pc_w913_buf           = pc_w913;


wire                             spc914_inst_done_buf  = spc914_inst_done;
wire [63:0]                      pc_w914_buf           = pc_w914;


wire                             spc915_inst_done_buf  = spc915_inst_done;
wire [63:0]                      pc_w915_buf           = pc_w915;


wire                             spc916_inst_done_buf  = spc916_inst_done;
wire [63:0]                      pc_w916_buf           = pc_w916;


wire                             spc917_inst_done_buf  = spc917_inst_done;
wire [63:0]                      pc_w917_buf           = pc_w917;


wire                             spc918_inst_done_buf  = spc918_inst_done;
wire [63:0]                      pc_w918_buf           = pc_w918;


wire                             spc919_inst_done_buf  = spc919_inst_done;
wire [63:0]                      pc_w919_buf           = pc_w919;


wire                             spc920_inst_done_buf  = spc920_inst_done;
wire [63:0]                      pc_w920_buf           = pc_w920;


wire                             spc921_inst_done_buf  = spc921_inst_done;
wire [63:0]                      pc_w921_buf           = pc_w921;


wire                             spc922_inst_done_buf  = spc922_inst_done;
wire [63:0]                      pc_w922_buf           = pc_w922;


wire                             spc923_inst_done_buf  = spc923_inst_done;
wire [63:0]                      pc_w923_buf           = pc_w923;


wire                             spc924_inst_done_buf  = spc924_inst_done;
wire [63:0]                      pc_w924_buf           = pc_w924;


wire                             spc925_inst_done_buf  = spc925_inst_done;
wire [63:0]                      pc_w925_buf           = pc_w925;


wire                             spc926_inst_done_buf  = spc926_inst_done;
wire [63:0]                      pc_w926_buf           = pc_w926;


wire                             spc927_inst_done_buf  = spc927_inst_done;
wire [63:0]                      pc_w927_buf           = pc_w927;


wire                             spc928_inst_done_buf  = spc928_inst_done;
wire [63:0]                      pc_w928_buf           = pc_w928;


wire                             spc929_inst_done_buf  = spc929_inst_done;
wire [63:0]                      pc_w929_buf           = pc_w929;


wire                             spc930_inst_done_buf  = spc930_inst_done;
wire [63:0]                      pc_w930_buf           = pc_w930;


wire                             spc931_inst_done_buf  = spc931_inst_done;
wire [63:0]                      pc_w931_buf           = pc_w931;


wire                             spc932_inst_done_buf  = spc932_inst_done;
wire [63:0]                      pc_w932_buf           = pc_w932;


wire                             spc933_inst_done_buf  = spc933_inst_done;
wire [63:0]                      pc_w933_buf           = pc_w933;


wire                             spc934_inst_done_buf  = spc934_inst_done;
wire [63:0]                      pc_w934_buf           = pc_w934;


wire                             spc935_inst_done_buf  = spc935_inst_done;
wire [63:0]                      pc_w935_buf           = pc_w935;


wire                             spc936_inst_done_buf  = spc936_inst_done;
wire [63:0]                      pc_w936_buf           = pc_w936;


wire                             spc937_inst_done_buf  = spc937_inst_done;
wire [63:0]                      pc_w937_buf           = pc_w937;


wire                             spc938_inst_done_buf  = spc938_inst_done;
wire [63:0]                      pc_w938_buf           = pc_w938;


wire                             spc939_inst_done_buf  = spc939_inst_done;
wire [63:0]                      pc_w939_buf           = pc_w939;


wire                             spc940_inst_done_buf  = spc940_inst_done;
wire [63:0]                      pc_w940_buf           = pc_w940;


wire                             spc941_inst_done_buf  = spc941_inst_done;
wire [63:0]                      pc_w941_buf           = pc_w941;


wire                             spc942_inst_done_buf  = spc942_inst_done;
wire [63:0]                      pc_w942_buf           = pc_w942;


wire                             spc943_inst_done_buf  = spc943_inst_done;
wire [63:0]                      pc_w943_buf           = pc_w943;


wire                             spc944_inst_done_buf  = spc944_inst_done;
wire [63:0]                      pc_w944_buf           = pc_w944;


wire                             spc945_inst_done_buf  = spc945_inst_done;
wire [63:0]                      pc_w945_buf           = pc_w945;


wire                             spc946_inst_done_buf  = spc946_inst_done;
wire [63:0]                      pc_w946_buf           = pc_w946;


wire                             spc947_inst_done_buf  = spc947_inst_done;
wire [63:0]                      pc_w947_buf           = pc_w947;


wire                             spc948_inst_done_buf  = spc948_inst_done;
wire [63:0]                      pc_w948_buf           = pc_w948;


wire                             spc949_inst_done_buf  = spc949_inst_done;
wire [63:0]                      pc_w949_buf           = pc_w949;


wire                             spc950_inst_done_buf  = spc950_inst_done;
wire [63:0]                      pc_w950_buf           = pc_w950;


wire                             spc951_inst_done_buf  = spc951_inst_done;
wire [63:0]                      pc_w951_buf           = pc_w951;


wire                             spc952_inst_done_buf  = spc952_inst_done;
wire [63:0]                      pc_w952_buf           = pc_w952;


wire                             spc953_inst_done_buf  = spc953_inst_done;
wire [63:0]                      pc_w953_buf           = pc_w953;


wire                             spc954_inst_done_buf  = spc954_inst_done;
wire [63:0]                      pc_w954_buf           = pc_w954;


wire                             spc955_inst_done_buf  = spc955_inst_done;
wire [63:0]                      pc_w955_buf           = pc_w955;


wire                             spc956_inst_done_buf  = spc956_inst_done;
wire [63:0]                      pc_w956_buf           = pc_w956;


wire                             spc957_inst_done_buf  = spc957_inst_done;
wire [63:0]                      pc_w957_buf           = pc_w957;


wire                             spc958_inst_done_buf  = spc958_inst_done;
wire [63:0]                      pc_w958_buf           = pc_w958;


wire                             spc959_inst_done_buf  = spc959_inst_done;
wire [63:0]                      pc_w959_buf           = pc_w959;


wire                             spc960_inst_done_buf  = spc960_inst_done;
wire [63:0]                      pc_w960_buf           = pc_w960;


wire                             spc961_inst_done_buf  = spc961_inst_done;
wire [63:0]                      pc_w961_buf           = pc_w961;


wire                             spc962_inst_done_buf  = spc962_inst_done;
wire [63:0]                      pc_w962_buf           = pc_w962;


wire                             spc963_inst_done_buf  = spc963_inst_done;
wire [63:0]                      pc_w963_buf           = pc_w963;


wire                             spc964_inst_done_buf  = spc964_inst_done;
wire [63:0]                      pc_w964_buf           = pc_w964;


wire                             spc965_inst_done_buf  = spc965_inst_done;
wire [63:0]                      pc_w965_buf           = pc_w965;


wire                             spc966_inst_done_buf  = spc966_inst_done;
wire [63:0]                      pc_w966_buf           = pc_w966;


wire                             spc967_inst_done_buf  = spc967_inst_done;
wire [63:0]                      pc_w967_buf           = pc_w967;


wire                             spc968_inst_done_buf  = spc968_inst_done;
wire [63:0]                      pc_w968_buf           = pc_w968;


wire                             spc969_inst_done_buf  = spc969_inst_done;
wire [63:0]                      pc_w969_buf           = pc_w969;


wire                             spc970_inst_done_buf  = spc970_inst_done;
wire [63:0]                      pc_w970_buf           = pc_w970;


wire                             spc971_inst_done_buf  = spc971_inst_done;
wire [63:0]                      pc_w971_buf           = pc_w971;


wire                             spc972_inst_done_buf  = spc972_inst_done;
wire [63:0]                      pc_w972_buf           = pc_w972;


wire                             spc973_inst_done_buf  = spc973_inst_done;
wire [63:0]                      pc_w973_buf           = pc_w973;


wire                             spc974_inst_done_buf  = spc974_inst_done;
wire [63:0]                      pc_w974_buf           = pc_w974;


wire                             spc975_inst_done_buf  = spc975_inst_done;
wire [63:0]                      pc_w975_buf           = pc_w975;


wire                             spc976_inst_done_buf  = spc976_inst_done;
wire [63:0]                      pc_w976_buf           = pc_w976;


wire                             spc977_inst_done_buf  = spc977_inst_done;
wire [63:0]                      pc_w977_buf           = pc_w977;


wire                             spc978_inst_done_buf  = spc978_inst_done;
wire [63:0]                      pc_w978_buf           = pc_w978;


wire                             spc979_inst_done_buf  = spc979_inst_done;
wire [63:0]                      pc_w979_buf           = pc_w979;


wire                             spc980_inst_done_buf  = spc980_inst_done;
wire [63:0]                      pc_w980_buf           = pc_w980;


wire                             spc981_inst_done_buf  = spc981_inst_done;
wire [63:0]                      pc_w981_buf           = pc_w981;


wire                             spc982_inst_done_buf  = spc982_inst_done;
wire [63:0]                      pc_w982_buf           = pc_w982;


wire                             spc983_inst_done_buf  = spc983_inst_done;
wire [63:0]                      pc_w983_buf           = pc_w983;


wire                             spc984_inst_done_buf  = spc984_inst_done;
wire [63:0]                      pc_w984_buf           = pc_w984;


wire                             spc985_inst_done_buf  = spc985_inst_done;
wire [63:0]                      pc_w985_buf           = pc_w985;


wire                             spc986_inst_done_buf  = spc986_inst_done;
wire [63:0]                      pc_w986_buf           = pc_w986;


wire                             spc987_inst_done_buf  = spc987_inst_done;
wire [63:0]                      pc_w987_buf           = pc_w987;


wire                             spc988_inst_done_buf  = spc988_inst_done;
wire [63:0]                      pc_w988_buf           = pc_w988;


wire                             spc989_inst_done_buf  = spc989_inst_done;
wire [63:0]                      pc_w989_buf           = pc_w989;


wire                             spc990_inst_done_buf  = spc990_inst_done;
wire [63:0]                      pc_w990_buf           = pc_w990;


wire                             spc991_inst_done_buf  = spc991_inst_done;
wire [63:0]                      pc_w991_buf           = pc_w991;


wire                             spc992_inst_done_buf  = spc992_inst_done;
wire [63:0]                      pc_w992_buf           = pc_w992;


wire                             spc993_inst_done_buf  = spc993_inst_done;
wire [63:0]                      pc_w993_buf           = pc_w993;


wire                             spc994_inst_done_buf  = spc994_inst_done;
wire [63:0]                      pc_w994_buf           = pc_w994;


wire                             spc995_inst_done_buf  = spc995_inst_done;
wire [63:0]                      pc_w995_buf           = pc_w995;


wire                             spc996_inst_done_buf  = spc996_inst_done;
wire [63:0]                      pc_w996_buf           = pc_w996;


wire                             spc997_inst_done_buf  = spc997_inst_done;
wire [63:0]                      pc_w997_buf           = pc_w997;


wire                             spc998_inst_done_buf  = spc998_inst_done;
wire [63:0]                      pc_w998_buf           = pc_w998;


wire                             spc999_inst_done_buf  = spc999_inst_done;
wire [63:0]                      pc_w999_buf           = pc_w999;


wire                             spc1000_inst_done_buf  = spc1000_inst_done;
wire [63:0]                      pc_w1000_buf           = pc_w1000;


wire                             spc1001_inst_done_buf  = spc1001_inst_done;
wire [63:0]                      pc_w1001_buf           = pc_w1001;


wire                             spc1002_inst_done_buf  = spc1002_inst_done;
wire [63:0]                      pc_w1002_buf           = pc_w1002;


wire                             spc1003_inst_done_buf  = spc1003_inst_done;
wire [63:0]                      pc_w1003_buf           = pc_w1003;


wire                             spc1004_inst_done_buf  = spc1004_inst_done;
wire [63:0]                      pc_w1004_buf           = pc_w1004;


wire                             spc1005_inst_done_buf  = spc1005_inst_done;
wire [63:0]                      pc_w1005_buf           = pc_w1005;


wire                             spc1006_inst_done_buf  = spc1006_inst_done;
wire [63:0]                      pc_w1006_buf           = pc_w1006;


wire                             spc1007_inst_done_buf  = spc1007_inst_done;
wire [63:0]                      pc_w1007_buf           = pc_w1007;


wire                             spc1008_inst_done_buf  = spc1008_inst_done;
wire [63:0]                      pc_w1008_buf           = pc_w1008;


wire                             spc1009_inst_done_buf  = spc1009_inst_done;
wire [63:0]                      pc_w1009_buf           = pc_w1009;


wire                             spc1010_inst_done_buf  = spc1010_inst_done;
wire [63:0]                      pc_w1010_buf           = pc_w1010;


wire                             spc1011_inst_done_buf  = spc1011_inst_done;
wire [63:0]                      pc_w1011_buf           = pc_w1011;


wire                             spc1012_inst_done_buf  = spc1012_inst_done;
wire [63:0]                      pc_w1012_buf           = pc_w1012;


wire                             spc1013_inst_done_buf  = spc1013_inst_done;
wire [63:0]                      pc_w1013_buf           = pc_w1013;


wire                             spc1014_inst_done_buf  = spc1014_inst_done;
wire [63:0]                      pc_w1014_buf           = pc_w1014;


wire                             spc1015_inst_done_buf  = spc1015_inst_done;
wire [63:0]                      pc_w1015_buf           = pc_w1015;


wire                             spc1016_inst_done_buf  = spc1016_inst_done;
wire [63:0]                      pc_w1016_buf           = pc_w1016;


wire                             spc1017_inst_done_buf  = spc1017_inst_done;
wire [63:0]                      pc_w1017_buf           = pc_w1017;


wire                             spc1018_inst_done_buf  = spc1018_inst_done;
wire [63:0]                      pc_w1018_buf           = pc_w1018;


wire                             spc1019_inst_done_buf  = spc1019_inst_done;
wire [63:0]                      pc_w1019_buf           = pc_w1019;


wire                             spc1020_inst_done_buf  = spc1020_inst_done;
wire [63:0]                      pc_w1020_buf           = pc_w1020;


wire                             spc1021_inst_done_buf  = spc1021_inst_done;
wire [63:0]                      pc_w1021_buf           = pc_w1021;


wire                             spc1022_inst_done_buf  = spc1022_inst_done;
wire [63:0]                      pc_w1022_buf           = pc_w1022;


wire                             spc1023_inst_done_buf  = spc1023_inst_done;
wire [63:0]                      pc_w1023_buf           = pc_w1023;




reg 	 ok_iob;
initial
begin
    ok_iob    = 0;
    fake_iob_out_data  = 0;
end

integer cpx_driven;

//// cmp clock domain
//// trin bug #65: use reference clock from the chip b/c the fake iob
//// needs to monitor the core PC
//always @(negedge `CHIP.clk_muxed)
//begin
//    if(ok_iob)
//    begin
            
//        cpx_driven = drive_iob();
//        if (cpx_driven) begin
//            fake_iob_out_data[`CPX_WIDTH-1:128] = get_cpx_word(0);
//            fake_iob_out_data[127:96] = get_cpx_word(1);
//            fake_iob_out_data[95:64] = get_cpx_word(2);
//            fake_iob_out_data[63:32] = get_cpx_word(3);
//            fake_iob_out_data[31:0] = get_cpx_word(4);
//            //$display("Doing IOB stuff - got values: %x %x %x %x %x", fake_iob_out_data[159:128], fake_iob_out_data[127:96], fake_iob_out_data[95:64], fake_iob_out_data[63:32], fake_iob_out_data[31:0]);
//        end else begin
//            fake_iob_out_data = {160{1'b0}};
//        end
//
//        // a little error check
//        if (iob_buffer_val && (out_buffer_val[out_write_index] | out_buffer_val[out_write_index + 1] == 1'b1))
//        begin
//            $display("%d : Simulation -> FAIL(%0s)", $time, "ciop_iob.v: IOB out buffer overflowed");
//            repeat(5)@(posedge clk);
//`ifndef DISABLE_ALL_MONITORS
//            `MONITOR_PATH.fail("ciop_iob.v: IOB out buffer overflowed");
//`endif
//        end
//    end // if (ok_iob)
//end // always @ (posedge cmp_gclk)

endmodule
