
import "DPI-C" function longint ColdDownThreshold_0_constantin_read();

module ColdDownThreshold_0_constantinReader(
  output reg [64 - 1:0] value
);

  initial value = ColdDownThreshold_0_constantin_read();
endmodule

import "DPI-C" function longint CorrectMissTrain0_constantin_read();

module CorrectMissTrain0_constantinReader(
  output reg [64 - 1:0] value
);

  initial value = CorrectMissTrain0_constantin_read();
endmodule

import "DPI-C" function longint depth0_constantin_read();

module depth0_constantinReader(
  output reg [64 - 1:0] value
);

  initial value = depth0_constantin_read();
endmodule

import "DPI-C" function longint enableDynamicPrefetcher0_constantin_read();

module enableDynamicPrefetcher0_constantinReader(
  output reg [64 - 1:0] value
);

  initial value = enableDynamicPrefetcher0_constantin_read();
endmodule

import "DPI-C" function longint ForceWriteLower_0_constantin_read();

module ForceWriteLower_0_constantinReader(
  output reg [64 - 1:0] value
);

  initial value = ForceWriteLower_0_constantin_read();
endmodule

import "DPI-C" function longint ForceWriteUpper_0_constantin_read();

module ForceWriteUpper_0_constantinReader(
  output reg [64 - 1:0] value
);

  initial value = ForceWriteUpper_0_constantin_read();
endmodule

import "DPI-C" function longint isFirstHitWrite0_constantin_read();

module isFirstHitWrite0_constantinReader(
  output reg [64 - 1:0] value
);

  initial value = isFirstHitWrite0_constantin_read();
endmodule

import "DPI-C" function longint isWriteBankConflictTable0_constantin_read();

module isWriteBankConflictTable0_constantinReader(
  output reg [64 - 1:0] value
);

  initial value = isWriteBankConflictTable0_constantin_read();
endmodule

import "DPI-C" function longint isWriteFetchToIBufferTable0_constantin_read();

module isWriteFetchToIBufferTable0_constantinReader(
  output reg [64 - 1:0] value
);

  initial value = isWriteFetchToIBufferTable0_constantin_read();
endmodule

import "DPI-C" function longint isWriteFTQTable0_constantin_read();

module isWriteFTQTable0_constantinReader(
  output reg [64 - 1:0] value
);

  initial value = isWriteFTQTable0_constantin_read();
endmodule

import "DPI-C" function longint isWriteICacheTable0_constantin_read();

module isWriteICacheTable0_constantinReader(
  output reg [64 - 1:0] value
);

  initial value = isWriteICacheTable0_constantin_read();
endmodule

import "DPI-C" function longint isWriteIfuWbToFtqTable0_constantin_read();

module isWriteIfuWbToFtqTable0_constantinReader(
  output reg [64 - 1:0] value
);

  initial value = isWriteIfuWbToFtqTable0_constantin_read();
endmodule

import "DPI-C" function longint isWriteInstInfoTable0_constantin_read();

module isWriteInstInfoTable0_constantinReader(
  output reg [64 - 1:0] value
);

  initial value = isWriteInstInfoTable0_constantin_read();
endmodule

import "DPI-C" function longint isWriteL1MissQMissTable0_constantin_read();

module isWriteL1MissQMissTable0_constantinReader(
  output reg [64 - 1:0] value
);

  initial value = isWriteL1MissQMissTable0_constantin_read();
endmodule

import "DPI-C" function longint isWriteL1TlbTable0_constantin_read();

module isWriteL1TlbTable0_constantinReader(
  output reg [64 - 1:0] value
);

  initial value = isWriteL1TlbTable0_constantin_read();
endmodule

import "DPI-C" function longint isWriteL2TlbMissQueueTable0_constantin_read();

module isWriteL2TlbMissQueueTable0_constantinReader(
  output reg [64 - 1:0] value
);

  initial value = isWriteL2TlbMissQueueTable0_constantin_read();
endmodule

import "DPI-C" function longint isWriteL2TlbPrefetchTable0_constantin_read();

module isWriteL2TlbPrefetchTable0_constantinReader(
  output reg [64 - 1:0] value
);

  initial value = isWriteL2TlbPrefetchTable0_constantin_read();
endmodule

import "DPI-C" function longint isWriteLoadAccessTable0_constantin_read();

module isWriteLoadAccessTable0_constantinReader(
  output reg [64 - 1:0] value
);

  initial value = isWriteLoadAccessTable0_constantin_read();
endmodule

import "DPI-C" function longint isWriteLoadMissTable0_constantin_read();

module isWriteLoadMissTable0_constantinReader(
  output reg [64 - 1:0] value
);

  initial value = isWriteLoadMissTable0_constantin_read();
endmodule

import "DPI-C" function longint isWritePageCacheTable0_constantin_read();

module isWritePageCacheTable0_constantinReader(
  output reg [64 - 1:0] value
);

  initial value = isWritePageCacheTable0_constantin_read();
endmodule

import "DPI-C" function longint isWritePrefetchPtrTable0_constantin_read();

module isWritePrefetchPtrTable0_constantinReader(
  output reg [64 - 1:0] value
);

  initial value = isWritePrefetchPtrTable0_constantin_read();
endmodule

import "DPI-C" function longint isWritePTWTable0_constantin_read();

module isWritePTWTable0_constantinReader(
  output reg [64 - 1:0] value
);

  initial value = isWritePTWTable0_constantin_read();
endmodule

import "DPI-C" function longint nMaxPrefetchEntry0_constantin_read();

module nMaxPrefetchEntry0_constantinReader(
  output reg [64 - 1:0] value
);

  initial value = nMaxPrefetchEntry0_constantin_read();
endmodule

import "DPI-C" function longint StoreBufferBase_0_constantin_read();

module StoreBufferBase_0_constantinReader(
  output reg [64 - 1:0] value
);

  initial value = StoreBufferBase_0_constantin_read();
endmodule

import "DPI-C" function longint StoreBufferThreshold_0_constantin_read();

module StoreBufferThreshold_0_constantinReader(
  output reg [64 - 1:0] value
);

  initial value = StoreBufferThreshold_0_constantin_read();
endmodule

import "DPI-C" function longint StoreWaitThreshold_0_constantin_read();

module StoreWaitThreshold_0_constantinReader(
  output reg [64 - 1:0] value
);

  initial value = StoreWaitThreshold_0_constantin_read();
endmodule
