/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module bootrom_linux (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [63:0]  addr_i,
   output logic [63:0]  rdata_o
);
    localparam int RomSize = 734;

    const logic [RomSize-1:0][63:0] mem = {
        64'h000000ff_f0c2c004,
        64'h000000ff_f0c2c003,
        64'h000000ff_f0c2c001,
        64'h000000ff_f0c2c005,
        64'h00000000_00000000,
        64'h0a0d2165_6e6f6420,
        64'h00000000_00206567,
        64'h616d6920_746f6f62,
        64'h20676e69_79706f63,
        64'h00000000_00000009,
        64'h3a656d61_6e090a0d,
        64'h00093a73_65747562,
        64'h69727474_61090a0d,
        64'h00000009_3a61626c,
        64'h20747361_6c090a0d,
        64'h0000093a_61626c20,
        64'h74737269_66090a0d,
        64'h00000000_00000000,
        64'h09202020_20203a64,
        64'h69756720_6e6f6974,
        64'h69747261_70090a0d,
        64'h00000000_00000000,
        64'h093a6469_75672065,
        64'h70797420_6e6f6974,
        64'h69747261_70090a0d,
        64'h00000000_20797274,
        64'h6e65206e_6f697469,
        64'h74726170_20747067,
        64'h00000009_20203a73,
        64'h65697274_6e65206e,
        64'h6f697469_74726170,
        64'h20657a69_73090a0d,
        64'h00000009_3a736569,
        64'h72746e65_206e6f69,
        64'h74697472_61702072,
        64'h65626d75_6e090a0d,
        64'h00000009_2020203a,
        64'h61626c20_73656972,
        64'h746e6520_6e6f6974,
        64'h69747261_70090a0d,
        64'h00093a61_646c2070,
        64'h756b6361_62090a0d,
        64'h00000000_00000000,
        64'h093a6162_6c20746e,
        64'h65727275_63090a0d,
        64'h00000009_3a646576,
        64'h72657365_72090a0d,
        64'h00093a72_65646165,
        64'h685f6372_63090a0d,
        64'h00000000_00000909,
        64'h3a657a69_73090a0d,
        64'h00000009_3a6e6f69,
        64'h73697665_72090a0d,
        64'h0000093a_65727574,
        64'h616e6769_73090a0d,
        64'h00000000_003a7265,
        64'h64616568_20656c62,
        64'h6174206e_6f697469,
        64'h74726170_20747067,
        64'h0000203a_65756c61,
        64'h76206e72_75746572,
        64'h2079706f_63206473,
        64'h00000000_0000000a,
        64'h0d216465_6c696166,
        64'h20647261_63204453,
        64'h00000000_0a0d676e,
        64'h69746978_65202e2e,
        64'h2e647320_657a696c,
        64'h61697469_6e692074,
        64'h6f6e2064_6c756f63,
        64'h00000000_00292520,
        64'h00000000_00000028,
        64'h20736b63_6f6c6220,
        64'h00000000_20666f20,
        64'h0000206b_636f6c62,
        64'h20676e69_79706f63,
        64'h00000000_00000008,
        64'h0000000a_0d202e2e,
        64'h2e445320_676e697a,
        64'h696c6169_74696e69,
        64'h00000000_203f3f79,
        64'h74706d65_20746f6e,
        64'h206f6669_66207872,
        64'h00000000_00000a0d,
        64'h2164657a_696c6169,
        64'h74696e69_20495053,
        64'h00000000_00007830,
        64'h203a7375_74617473,
        64'h00000000_00000a0d,
        64'h49505320_74696e69,
        64'h00000000_0000000a,
        64'h0d216465_7a696c61,
        64'h6974696e_69206473,
        64'h00000000_00007665,
        64'h646e2c76_63736972,
        64'h00797469_726f6972,
        64'h702d7861_6d2c7663,
        64'h73697200_73656d61,
        64'h6e2d6765_72006465,
        64'h646e6574_78652d73,
        64'h74707572_7265746e,
        64'h69007466_6968732d,
        64'h67657200_73747075,
        64'h72726574_6e690074,
        64'h6e657261_702d7470,
        64'h75727265_746e6900,
        64'h64656570_732d746e,
        64'h65727275_6300656c,
        64'h646e6168_70007265,
        64'h6c6c6f72_746e6f63,
        64'h2d747075_72726574,
        64'h6e690073_6c6c6563,
        64'h2d747075_72726574,
        64'h6e692300_74696c70,
        64'h732d626c_74006570,
        64'h79742d75_6d6d0061,
        64'h73692c76_63736972,
        64'h00737574_61747300,
        64'h67657200_65707974,
        64'h5f656369_76656400,
        64'h79636e65_75716572,
        64'h662d6b63_6f6c6300,
        64'h79636e65_75716572,
        64'h662d6573_6162656d,
        64'h69740030_6c616972,
        64'h65730065_6c6f736e,
        64'h6f630068_7461702d,
        64'h74756f64_74730065,
        64'h6c626974_61706d6f,
        64'h6300636f_6c65722d,
        64'h6572702d_6d642c74,
        64'h6f6f622d_7500736c,
        64'h6c65632d_657a6973,
        64'h2300736c_6c65632d,
        64'h73736572_64646123,
        64'h09000000_02000000,
        64'h02000000_01000000,
        64'hd3000000_04000000,
        64'h03000000_01000000,
        64'h40010000_04000000,
        64'h03000000_07000000,
        64'h2d010000_04000000,
        64'h03000000_00000004,
        64'h00000000_000010f1,
        64'hff000000_85000000,
        64'h10000000_03000000,
        64'h09000000_02000000,
        64'h0b000000_02000000,
        64'h0f010000_10000000,
        64'h03000000_be000000,
        64'h00000000_03000000,
        64'h00306369_6c702c76,
        64'h63736972_2f000000,
        64'h0c000000_03000000,
        64'h01000000_ad000000,
        64'h04000000_03000000,
        64'h00000000_00000000,
        64'h04000000_03000000,
        64'h1b000000_00000000,
        64'h03000000_00303030,
        64'h30303131_66666640,
        64'h63696c70_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_23010000,
        64'h08000000_03000000,
        64'h00000c00_00000000,
        64'h000002f1_ff000000,
        64'h85000000_10000000,
        64'h03000000_07000000,
        64'h02000000_03000000,
        64'h02000000_0f010000,
        64'h10000000_03000000,
        64'h00000000_30746e69,
        64'h6c632c76_63736972,
        64'h2f000000_0d000000,
        64'h03000000_1b000000,
        64'h00000000_03000000,
        64'h00000000_30303030,
        64'h32303166_66664074,
        64'h6e696c63_01000000,
        64'h02000000_00000000,
        64'h05010000_04000000,
        64'h03000000_01000000,
        64'hfa000000_04000000,
        64'h03000000_01000000,
        64'he9000000_04000000,
        64'h03000000_00c20100,
        64'hdb000000_04000000,
        64'h03000000_80f0fa02,
        64'h69000000_04000000,
        64'h03000000_00400d00,
        64'h00000000_00c0c2f0,
        64'hff000000_85000000,
        64'h10000000_03000000,
        64'h00303535_3631736e,
        64'h2f000000_08000000,
        64'h03000000_1b000000,
        64'h00000000_03000000,
        64'h00303030_63326330,
        64'h66666640_74726175,
        64'h01000000_02000000,
        64'h00000040_00000000,
        64'h00000080_00000000,
        64'h85000000_10000000,
        64'h03000000_00007972,
        64'h6f6d656d_79000000,
        64'h07000000_03000000,
        64'h1b000000_00000000,
        64'h03000000_00303030,
        64'h30303030_38407972,
        64'h6f6d656d_01000000,
        64'h02000000_02000000,
        64'h02000000_02000000,
        64'hd3000000_04000000,
        64'h03000000_00006374,
        64'h6e692d75_70632c76,
        64'h63736972_2f000000,
        64'h0f000000_03000000,
        64'hbe000000_00000000,
        64'h03000000_01000000,
        64'had000000_04000000,
        64'h03000000_00000000,
        64'h72656c6c_6f72746e,
        64'h6f632d74_70757272,
        64'h65746e69_01000000,
        64'ha3000000_00000000,
        64'h03000000_00003933,
        64'h76732c76_63736972,
        64'h9a000000_0b000000,
        64'h03000000_00006364,
        64'h66616d69_34367672,
        64'h90000000_0b000000,
        64'h03000000_00766373,
        64'h69720036_61766320,
        64'h2c70756f_72677768,
        64'h6e65706f_2f000000,
        64'h18000000_03000000,
        64'h00000000_79616b6f,
        64'h89000000_05000000,
        64'h03000000_00000000,
        64'h85000000_04000000,
        64'h03000000_00757063,
        64'h79000000_04000000,
        64'h03000000_1b000000,
        64'h00000000_03000000,
        64'h80f0fa02_69000000,
        64'h04000000_03000000,
        64'h00000030_40757063,
        64'h01000000_e1f50500,
        64'h56000000_04000000,
        64'h03000000_1b000000,
        64'h00000000_03000000,
        64'h00000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00000000_73757063,
        64'h01000000_02000000,
        64'h00000000_30303063,
        64'h32633066_66664074,
        64'h7261752f_4e000000,
        64'h11000000_03000000,
        64'h00000000_30303063,
        64'h32633066_66664074,
        64'h7261752f_46000000,
        64'h11000000_03000000,
        64'h1b000000_00000000,
        64'h03000000_00736573,
        64'h61696c61_01000000,
        64'h02000000_00000000,
        64'h30303235_31313a30,
        64'h74726175_3a000000,
        64'h0d000000_03000000,
        64'h1b000000_00000000,
        64'h03000000_00006e65,
        64'h736f6863_01000000,
        64'h00006d72_6f667461,
        64'h6c703661_76632c6e,
        64'h6f746970_6e65706f,
        64'h2f000000_17000000,
        64'h03000000_1b000000,
        64'h00000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00000000_01000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'hc0040000_4b010000,
        64'h00000000_10000000,
        64'h11000000_28000000,
        64'hf8040000_38000000,
        64'h43060000_edfe0dd0,
        64'h00000000_00000000,
        64'h00000000_00000a0d,
        64'h0a0d0a0d_2d2d2d2d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h2d2d2d2d_0a0d2020,
        64'h20202020_20202020,
        64'h34202f20_426b2034,
        64'h36202020_3a636f73,
        64'h7341202f_20657a69,
        64'h53202032_4c0a0d20,
        64'h20202020_20202020,
        64'h2034202f_20426b20,
        64'h38202020_203a636f,
        64'h73734120_2f20657a,
        64'h69532035_314c0a0d,
        64'h20202020_20202020,
        64'h20203420_2f20426b,
        64'h20382020_20203a63,
        64'h6f737341_202f2065,
        64'h7a695320_44314c0a,
        64'h0d202020_20202020,
        64'h20202034_202f2042,
        64'h6b203631_2020203a,
        64'h636f7373_41202f20,
        64'h657a6953_2049314c,
        64'h0a0d2020_20202020,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h20200a0d_20202020,
        64'h20202020_20202020,
        64'h20202020_424d2034,
        64'h32303120_20202020,
        64'h20202020_3a657a69,
        64'h53204d41_52440a0d,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h20202068_73656d5f,
        64'h64322020_20202020,
        64'h20202020_203a6b72,
        64'h6f777465_4e0a0d20,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h20206e77_6f6e6b6e,
        64'h55202020_20202020,
        64'h20203a71_65724620,
        64'h65726f43_0a0d2020,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h20312020_20202020,
        64'h20202020_20203a73,
        64'h65726f43_230a0d20,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h20203120_20202020,
        64'h20202020_203a7365,
        64'h6c69542d_59230a0d,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h20202031_20202020,
        64'h20202020_20203a73,
        64'h656c6954_2d58230a,
        64'h0d202020_20202020,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h200a0d20_20202020,
        64'h20202020_20202020,
        64'h20202020_20203435,
        64'h3a34313a_33312035,
        64'h32303220_32312072,
        64'h614d2020_20202020,
        64'h20203a65_74614420,
        64'h646c6975_420a0d20,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h2020296e_6f697461,
        64'h6c756d69_53282065,
        64'h6e6f4e20_20202020,
        64'h2020203a_6472616f,
        64'h42204147_50460a0d,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h0a0d2020_20202020,
        64'h20202020_20202020,
        64'h20202020_20273461,
        64'h35356137_63322762,
        64'h20202020_3a6e6f69,
        64'h73726556_20656e61,
        64'h6972410a_0d202020,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h27396133_62366165,
        64'h30276220_3a6e6f69,
        64'h73726556_206e6f74,
        64'h69506e65_704f0a0d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h0a0d2d2d_20202020,
        64'h20206d72_6f667461,
        64'h6c502065_6e616972,
        64'h412b6e6f_7469506e,
        64'h65704f20_20202020,
        64'h2d2d0a0d_2d2d2d2d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h2d2d2d2d_0a0d0a0d,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h46454443_42413938,
        64'h37363534_33323130,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_80820141,
        64'h450160a2_cfdff0ef,
        64'h057e65c1_45058ebf,
        64'hf0efb5a5_05130000,
        64'h15178f7f_f0ef15e5,
        64'h05130000_05178a9f,
        64'hf0efe406_38050513,
        64'h20058593_114101c9,
        64'hc53765f1_b39591bf,
        64'hf0efe425_05130000,
        64'h1517bbd9_bdc50513,
        64'h00001517_a3dff0ef,
        64'h854a937f_f0efc9e5,
        64'h05130000_1517943f,
        64'hf0efc925_05130000,
        64'h1517bbfd_c0450513,
        64'h00001517_a65ff0ef,
        64'h852695ff_f0efcc65,
        64'h05130000_151796bf,
        64'hf0efcba5_05130000,
        64'h1517c929_84aac97f,
        64'hf0ef8552_8656020b,
        64'h2583987f_f0efc3e5,
        64'h05130000_1517993f,
        64'hf0efea25_05130000,
        64'h1517f579_10e30804,
        64'h84939a7f_f0ef2905,
        64'hc6050513_00001517,
        64'hff999be3_b09ff0ef,
        64'h09850009_c5039c3f,
        64'hf0efec25_05130000,
        64'h1517adbf_f0ef6888,
        64'h9d5ff0ef_ec450513,
        64'h00001517_aedff0ef,
        64'h64889e7f_f0efec65,
        64'h05130000_1517afff,
        64'hf0ef0604_8c930184,
        64'h89936088_a01ff0ef,
        64'hed050513_00001517,
        64'hfe999be3_b61ff0ef,
        64'h09850009_c503ff04,
        64'h8993a1ff_f0efece5,
        64'h05130000_1517ff89,
        64'h99e3b7ff_f0ef0985,
        64'h0007c503_013c87b3,
        64'h4981a3ff_f0effe04,
        64'h8c93ed25_05130000,
        64'h1517b9ff_f0ef0ff9,
        64'h7513a57f_f0efece5,
        64'h05130000_15174b91,
        64'h4c411005_1e631004,
        64'h892a8b0a_d8dff0ef,
        64'h850a4605_71010489,
        64'h2583a7ff_f0efd365,
        64'h05130000_1517b55f,
        64'hf0ef4556_a91ff0ef,
        64'hee850513_00001517,
        64'hb67ff0ef_4546aa3f,
        64'hf0efeda5_05130000,
        64'h1517bbbf_f0ef6526,
        64'hab5ff0ef_ecc50513,
        64'h00001517_bcdff0ef,
        64'h7502ac7f_f0efece5,
        64'h05130000_1517bdff,
        64'hf0ef6562_ad9ff0ef,
        64'hec850513_00001517,
        64'hbafff0ef_4552aebf,
        64'hf0efeca5_05130000,
        64'h1517bc1f_f0ef4542,
        64'hafdff0ef_ecc50513,
        64'h00001517_bd3ff0ef,
        64'h4532b0ff_f0efece5,
        64'h05130000_1517be5f,
        64'hf0ef4522_b21ff0ef,
        64'hed050513_00001517,
        64'hc39ff0ef_6502b33f,
        64'hf0efed25_05130000,
        64'h1517b3ff_f0efebe5,
        64'h05130000_1517bf59,
        64'h54f9b4ff_f0efe065,
        64'h05130000_1517c67f,
        64'hf0ef8526_b61ff0ef,
        64'hec850513_00001517,
        64'hb6dff0ef_ebc50513,
        64'h00001517_c90584aa,
        64'h890ae9bf_f0ef850a,
        64'h45854605_7101b8bf,
        64'hf0efdfa5_05130000,
        64'h15178082_61256ca2,
        64'h6c426be2_7b027aa2,
        64'h7a4279e2_690664a6,
        64'h64468526_60e6fa04,
        64'h011354fd_bb9ff0ef,
        64'hee050513_00001517,
        64'hc905ecbf_f0ef8aae,
        64'h8a2a1080_e466e862,
        64'hec5ef05a_fc4ee0ca,
        64'he4a6ec86_f456f852,
        64'he8a2711d_b7bd2c05,
        64'hbedff0ef_edc50513,
        64'h00001517_b7a10b85,
        64'h20048493_ff5799e3,
        64'he29007a1_00e786b3,
        64'h621000f4_86334781,
        64'h974e009b_97139c29,
        64'hc1dff0ef_f3c50513,
        64'h00001517_9c29c7df,
        64'hf0ef0325_553b4585,
        64'h036a053b_9c29c3bf,
        64'hf0eff4a5_05130000,
        64'h15179c29_c9bff0ef,
        64'h854a9c29_4585c53f,
        64'hf0eff5a5_05130000,
        64'h15179c29_cb3ff0ef,
        64'h855a0005_041b4585,
        64'hc6dff0ef_f6450513,
        64'h00001517_09841263,
        64'h060c1363_034b7c3b,
        64'h80826161_45016c02,
        64'h6ba26b42_6ae27a02,
        64'h79a27942_74e26406,
        64'h60a6c9ff_f0eff565,
        64'h05130000_1517032b,
        64'h6563000b_8b1b2000,
        64'h0a930640_0a134401,
        64'h4b8100f5_84b38932,
        64'h89aae062_e85ae486,
        64'he45eec56_f052f44e,
        64'hf84afc26_e0a21792,
        64'h715d47bd_0177d593,
        64'h02059793_80820141,
        64'h450160a2_cf1ff0ef,
        64'he406fcc5_05131141,
        64'h00001517_8082557d,
        64'hb7d900d7_00230785,
        64'h00f60733_06c82683,
        64'hff698b05_5178b77d,
        64'hd6b80785_00074703,
        64'h00f50733_80824501,
        64'hd3b84719_dbb8577d,
        64'h200007b7_02b6e163,
        64'h0007869b_20000837,
        64'h20000537_fff58b85,
        64'h537c2000_0737d3b8,
        64'h200007b7_10600713,
        64'hfff537fd_00010320,
        64'h079304b7_61630007,
        64'h871b4781_200006b7,
        64'hdbb85779_200007b7,
        64'h06b7ee63_10000793,
        64'h80826105_64a2d3b8,
        64'h4719dbb8_64420ff4,
        64'h7513577d_200007b7,
        64'h60e2d9ff_f0ef0565,
        64'h05130000_1517eb7f,
        64'hf0ef9101_15024088,
        64'hdb5ff0ef_07450513,
        64'h00001517_e3958b85,
        64'h53fc57e0_ff658b05,
        64'h06478493_53f8d3b8,
        64'h10600713_200007b7,
        64'hfff537fd_00010640,
        64'h0793d7a8_dbb85779,
        64'he426e822_ec062000,
        64'h07b71101_bbdd6105,
        64'h0a050513_00001517,
        64'h64a260e2_6442d03c,
        64'h4799e0ff_f0ef0c65,
        64'h05130000_1517f27f,
        64'hf0ef9101_02049513,
        64'he25ff0ef_0bc50513,
        64'h00001517_5064d03c,
        64'h16600793_e39ff0ef,
        64'h0f050513_00001517,
        64'hf51ff0ef_91010204,
        64'h9513e4ff_f0ef0e65,
        64'h05130000_15175064,
        64'hd03c1040_07932000,
        64'h0437fff5_37fd0001,
        64'h47a9c3b8_47292000,
        64'h07b7e77f_f0efe426,
        64'he822ec06_10650513,
        64'h11010000_15178082,
        64'h41088082_c10c8082,
        64'h61054509_60e2e1ff,
        64'hf0ef0091_4503e27f,
        64'hf0ef0081_4503ed9f,
        64'hf0efec06_002c1101,
        64'h80826145_45416942,
        64'h64e27402_70a2ff24,
        64'h10e3e4bf_f0ef0091,
        64'h4503e53f_f0ef3461,
        64'h00814503_f07ff0ef,
        64'h0ff57513_002c0084,
        64'hd5335961_03800413,
        64'h84aaf406_e84aec26,
        64'hf0227179_80826145,
        64'h45216942_64e27402,
        64'h70a2ff24_10e3e8ff,
        64'hf0ef0091_4503e97f,
        64'hf0ef3461_00814503,
        64'hf4bff0ef_0ff57513,
        64'h002c0084_d53b5961,
        64'h446184aa_f406e84a,
        64'hec26f022_71798082,
        64'h612169e2_854e6b02,
        64'h6aa26a42_790274a2,
        64'h744270e2_fd5913e3,
        64'h397d85d2_eddff0ef,
        64'h0007c503_97ba8bbd,
        64'h02d7d7bb_29856ce7,
        64'h07130000_071702ba,
        64'h706300d7_f4630364,
        64'h543b0009_0a1b0284,
        64'hf4bb0004_069b0004,
        64'h879b5afd_4b294981,
        64'h4925a004_041384aa,
        64'he852fc06_e05ae456,
        64'hec4ef04a_f4263b9a,
        64'hd437f822_71398082,
        64'h00f58023_0007c783,
        64'h00e580a3_97aa8111,
        64'h00074703_973e00f5,
        64'h77137327_87930000,
        64'h0797b7c5_f5dff0ef,
        64'h853e8082_610564a2,
        64'h644260e2_e791fff7,
        64'hc7830084_87b30405,
        64'h0004051b_440184aa,
        64'hec06e426_e8221101,
        64'h808200e7_80230200,
        64'h071355a7_b7830000,
        64'h179700f7_0023478d,
        64'h00a68023_0ff57513,
        64'h00c78023_0085551b,
        64'h0ff57613_07ba30b7,
        64'h879303ff_c7b700f7,
        64'h0023f800_07930006,
        64'h802358a7_b7030000,
        64'h179758a7_b6830000,
        64'h179702b5_553b0045,
        64'h959b8082_00a78023,
        64'h07ba30b7_879303ff,
        64'hc7b7dbe5_0207f793,
        64'h0007c783_5ac7b783,
        64'h00001797_80820205,
        64'h75130007_c5035be7,
        64'hb7830000_17978082,
        64'h0ff57513_00054503,
        64'h808200b5_00238082,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00048067_01f49493,
        64'h0010049b_d5c58593,
        64'h00001597_f1402573,
        64'hff2496e3_00100493,
        64'h0004a903_04048493,
        64'h01a49493_0210049b,
        64'h0924a4af_00090913,
        64'h00190913_04048493,
        64'h01a49493_0210049b,
        64'hff2496e3_f14024f3,
        64'h0004a903_04048493,
        64'h01a49493_0210049b,
        64'h079000ef_01a11113,
        64'h0210011b_01249863,
        64'hf1402973_00000493
    };

    logic [$clog2(RomSize)-1:0] addr_q;

    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
        end
    end

    // this prevents spurious Xes from propagating into
    // the speculative fetch stage of the core
    assign rdata_o = (addr_q < RomSize) ? mem[addr_q] : '0;
endmodule
