// Modified by Princeton University on June 9th, 2015
// ========== Copyright Header Begin ==========================================
//
// OpenSPARC T1 Processor File: pc_cmp.v
// Copyright (c) 2006 Sun Microsystems, Inc.  All Rights Reserved.
// DO NOT ALTER OR REMOVE COPYRIGHT NOTICES.
//
// The above named program is free software; you can redistribute it and/or
// modify it under the terms of the GNU General Public
// License version 2 as published by the Free Software Foundation.
//
// The above named program is distributed in the hope that it will be
// useful, but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
// General Public License for more details.
//
// You should have received a copy of the GNU General Public
// License along with this work; if not, write to the Free Software
// Foundation, Inc., 51 Franklin St, Fifth Floor, Boston, MA 02110-1301, USA.
//
// ========== Copyright Header End ============================================

`include "define.tmp.h"
`include "ifu.tmp.h"

// /home/gl/work/openpiton/piton/verif/env/manycore/devices_ariane.xml
`define GOOD_TRAP_COUNTER 1


 module pc_cmp(/*AUTOARG*/
     // Inputs
     clk,
     rst_l
 );
input clk;
input rst_l;

// trap register

reg [4095:0]   active_thread;
reg [4:0]    thread_status[4095:0];

reg [1023:0]   good = '0;
reg [1023:0]   done;

reg [31:0]     timeout [4095:0];


reg [63:0]    good_trap[`GOOD_TRAP_COUNTER-1:0];
reg [63:0]    bad_trap [`GOOD_TRAP_COUNTER-1:0];

reg [`GOOD_TRAP_COUNTER-1:0] good_trap_exists;
reg [`GOOD_TRAP_COUNTER-1:0] bad_trap_exists;

reg           dum;
reg           hit_bad = 0;

integer       time_tmp, trap_count;


    reg spc0_inst_done;
    wire [1:0]   spc0_thread_id;
    wire [63:0]      spc0_rtl_pc;
    wire sas_m0;
    reg [63:0] spc0_phy_pc_w;

    

    reg spc1_inst_done;
    wire [1:0]   spc1_thread_id;
    wire [63:0]      spc1_rtl_pc;
    wire sas_m1;
    reg [63:0] spc1_phy_pc_w;

    

    reg spc2_inst_done;
    wire [1:0]   spc2_thread_id;
    wire [63:0]      spc2_rtl_pc;
    wire sas_m2;
    reg [63:0] spc2_phy_pc_w;

    

    reg spc3_inst_done;
    wire [1:0]   spc3_thread_id;
    wire [63:0]      spc3_rtl_pc;
    wire sas_m3;
    reg [63:0] spc3_phy_pc_w;

    

    reg spc4_inst_done;
    wire [1:0]   spc4_thread_id;
    wire [63:0]      spc4_rtl_pc;
    wire sas_m4;
    reg [63:0] spc4_phy_pc_w;

    

    reg spc5_inst_done;
    wire [1:0]   spc5_thread_id;
    wire [63:0]      spc5_rtl_pc;
    wire sas_m5;
    reg [63:0] spc5_phy_pc_w;

    

    reg spc6_inst_done;
    wire [1:0]   spc6_thread_id;
    wire [63:0]      spc6_rtl_pc;
    wire sas_m6;
    reg [63:0] spc6_phy_pc_w;

    

    reg spc7_inst_done;
    wire [1:0]   spc7_thread_id;
    wire [63:0]      spc7_rtl_pc;
    wire sas_m7;
    reg [63:0] spc7_phy_pc_w;

    

    reg spc8_inst_done;
    wire [1:0]   spc8_thread_id;
    wire [63:0]      spc8_rtl_pc;
    wire sas_m8;
    reg [63:0] spc8_phy_pc_w;

    

    reg spc9_inst_done;
    wire [1:0]   spc9_thread_id;
    wire [63:0]      spc9_rtl_pc;
    wire sas_m9;
    reg [63:0] spc9_phy_pc_w;

    

    reg spc10_inst_done;
    wire [1:0]   spc10_thread_id;
    wire [63:0]      spc10_rtl_pc;
    wire sas_m10;
    reg [63:0] spc10_phy_pc_w;

    

    reg spc11_inst_done;
    wire [1:0]   spc11_thread_id;
    wire [63:0]      spc11_rtl_pc;
    wire sas_m11;
    reg [63:0] spc11_phy_pc_w;

    

    reg spc12_inst_done;
    wire [1:0]   spc12_thread_id;
    wire [63:0]      spc12_rtl_pc;
    wire sas_m12;
    reg [63:0] spc12_phy_pc_w;

    

    reg spc13_inst_done;
    wire [1:0]   spc13_thread_id;
    wire [63:0]      spc13_rtl_pc;
    wire sas_m13;
    reg [63:0] spc13_phy_pc_w;

    

    reg spc14_inst_done;
    wire [1:0]   spc14_thread_id;
    wire [63:0]      spc14_rtl_pc;
    wire sas_m14;
    reg [63:0] spc14_phy_pc_w;

    

    reg spc15_inst_done;
    wire [1:0]   spc15_thread_id;
    wire [63:0]      spc15_rtl_pc;
    wire sas_m15;
    reg [63:0] spc15_phy_pc_w;

    

    reg spc16_inst_done;
    wire [1:0]   spc16_thread_id;
    wire [63:0]      spc16_rtl_pc;
    wire sas_m16;
    reg [63:0] spc16_phy_pc_w;

    

    reg spc17_inst_done;
    wire [1:0]   spc17_thread_id;
    wire [63:0]      spc17_rtl_pc;
    wire sas_m17;
    reg [63:0] spc17_phy_pc_w;

    

    reg spc18_inst_done;
    wire [1:0]   spc18_thread_id;
    wire [63:0]      spc18_rtl_pc;
    wire sas_m18;
    reg [63:0] spc18_phy_pc_w;

    

    reg spc19_inst_done;
    wire [1:0]   spc19_thread_id;
    wire [63:0]      spc19_rtl_pc;
    wire sas_m19;
    reg [63:0] spc19_phy_pc_w;

    

    reg spc20_inst_done;
    wire [1:0]   spc20_thread_id;
    wire [63:0]      spc20_rtl_pc;
    wire sas_m20;
    reg [63:0] spc20_phy_pc_w;

    

    reg spc21_inst_done;
    wire [1:0]   spc21_thread_id;
    wire [63:0]      spc21_rtl_pc;
    wire sas_m21;
    reg [63:0] spc21_phy_pc_w;

    

    reg spc22_inst_done;
    wire [1:0]   spc22_thread_id;
    wire [63:0]      spc22_rtl_pc;
    wire sas_m22;
    reg [63:0] spc22_phy_pc_w;

    

    reg spc23_inst_done;
    wire [1:0]   spc23_thread_id;
    wire [63:0]      spc23_rtl_pc;
    wire sas_m23;
    reg [63:0] spc23_phy_pc_w;

    

    reg spc24_inst_done;
    wire [1:0]   spc24_thread_id;
    wire [63:0]      spc24_rtl_pc;
    wire sas_m24;
    reg [63:0] spc24_phy_pc_w;

    

    reg spc25_inst_done;
    wire [1:0]   spc25_thread_id;
    wire [63:0]      spc25_rtl_pc;
    wire sas_m25;
    reg [63:0] spc25_phy_pc_w;

    

    reg spc26_inst_done;
    wire [1:0]   spc26_thread_id;
    wire [63:0]      spc26_rtl_pc;
    wire sas_m26;
    reg [63:0] spc26_phy_pc_w;

    

    reg spc27_inst_done;
    wire [1:0]   spc27_thread_id;
    wire [63:0]      spc27_rtl_pc;
    wire sas_m27;
    reg [63:0] spc27_phy_pc_w;

    

    reg spc28_inst_done;
    wire [1:0]   spc28_thread_id;
    wire [63:0]      spc28_rtl_pc;
    wire sas_m28;
    reg [63:0] spc28_phy_pc_w;

    

    reg spc29_inst_done;
    wire [1:0]   spc29_thread_id;
    wire [63:0]      spc29_rtl_pc;
    wire sas_m29;
    reg [63:0] spc29_phy_pc_w;

    

    reg spc30_inst_done;
    wire [1:0]   spc30_thread_id;
    wire [63:0]      spc30_rtl_pc;
    wire sas_m30;
    reg [63:0] spc30_phy_pc_w;

    

    reg spc31_inst_done;
    wire [1:0]   spc31_thread_id;
    wire [63:0]      spc31_rtl_pc;
    wire sas_m31;
    reg [63:0] spc31_phy_pc_w;

    

    reg spc32_inst_done;
    wire [1:0]   spc32_thread_id;
    wire [63:0]      spc32_rtl_pc;
    wire sas_m32;
    reg [63:0] spc32_phy_pc_w;

    

    reg spc33_inst_done;
    wire [1:0]   spc33_thread_id;
    wire [63:0]      spc33_rtl_pc;
    wire sas_m33;
    reg [63:0] spc33_phy_pc_w;

    

    reg spc34_inst_done;
    wire [1:0]   spc34_thread_id;
    wire [63:0]      spc34_rtl_pc;
    wire sas_m34;
    reg [63:0] spc34_phy_pc_w;

    

    reg spc35_inst_done;
    wire [1:0]   spc35_thread_id;
    wire [63:0]      spc35_rtl_pc;
    wire sas_m35;
    reg [63:0] spc35_phy_pc_w;

    

    reg spc36_inst_done;
    wire [1:0]   spc36_thread_id;
    wire [63:0]      spc36_rtl_pc;
    wire sas_m36;
    reg [63:0] spc36_phy_pc_w;

    

    reg spc37_inst_done;
    wire [1:0]   spc37_thread_id;
    wire [63:0]      spc37_rtl_pc;
    wire sas_m37;
    reg [63:0] spc37_phy_pc_w;

    

    reg spc38_inst_done;
    wire [1:0]   spc38_thread_id;
    wire [63:0]      spc38_rtl_pc;
    wire sas_m38;
    reg [63:0] spc38_phy_pc_w;

    

    reg spc39_inst_done;
    wire [1:0]   spc39_thread_id;
    wire [63:0]      spc39_rtl_pc;
    wire sas_m39;
    reg [63:0] spc39_phy_pc_w;

    

    reg spc40_inst_done;
    wire [1:0]   spc40_thread_id;
    wire [63:0]      spc40_rtl_pc;
    wire sas_m40;
    reg [63:0] spc40_phy_pc_w;

    

    reg spc41_inst_done;
    wire [1:0]   spc41_thread_id;
    wire [63:0]      spc41_rtl_pc;
    wire sas_m41;
    reg [63:0] spc41_phy_pc_w;

    

    reg spc42_inst_done;
    wire [1:0]   spc42_thread_id;
    wire [63:0]      spc42_rtl_pc;
    wire sas_m42;
    reg [63:0] spc42_phy_pc_w;

    

    reg spc43_inst_done;
    wire [1:0]   spc43_thread_id;
    wire [63:0]      spc43_rtl_pc;
    wire sas_m43;
    reg [63:0] spc43_phy_pc_w;

    

    reg spc44_inst_done;
    wire [1:0]   spc44_thread_id;
    wire [63:0]      spc44_rtl_pc;
    wire sas_m44;
    reg [63:0] spc44_phy_pc_w;

    

    reg spc45_inst_done;
    wire [1:0]   spc45_thread_id;
    wire [63:0]      spc45_rtl_pc;
    wire sas_m45;
    reg [63:0] spc45_phy_pc_w;

    

    reg spc46_inst_done;
    wire [1:0]   spc46_thread_id;
    wire [63:0]      spc46_rtl_pc;
    wire sas_m46;
    reg [63:0] spc46_phy_pc_w;

    

    reg spc47_inst_done;
    wire [1:0]   spc47_thread_id;
    wire [63:0]      spc47_rtl_pc;
    wire sas_m47;
    reg [63:0] spc47_phy_pc_w;

    

    reg spc48_inst_done;
    wire [1:0]   spc48_thread_id;
    wire [63:0]      spc48_rtl_pc;
    wire sas_m48;
    reg [63:0] spc48_phy_pc_w;

    

    reg spc49_inst_done;
    wire [1:0]   spc49_thread_id;
    wire [63:0]      spc49_rtl_pc;
    wire sas_m49;
    reg [63:0] spc49_phy_pc_w;

    

    reg spc50_inst_done;
    wire [1:0]   spc50_thread_id;
    wire [63:0]      spc50_rtl_pc;
    wire sas_m50;
    reg [63:0] spc50_phy_pc_w;

    

    reg spc51_inst_done;
    wire [1:0]   spc51_thread_id;
    wire [63:0]      spc51_rtl_pc;
    wire sas_m51;
    reg [63:0] spc51_phy_pc_w;

    

    reg spc52_inst_done;
    wire [1:0]   spc52_thread_id;
    wire [63:0]      spc52_rtl_pc;
    wire sas_m52;
    reg [63:0] spc52_phy_pc_w;

    

    reg spc53_inst_done;
    wire [1:0]   spc53_thread_id;
    wire [63:0]      spc53_rtl_pc;
    wire sas_m53;
    reg [63:0] spc53_phy_pc_w;

    

    reg spc54_inst_done;
    wire [1:0]   spc54_thread_id;
    wire [63:0]      spc54_rtl_pc;
    wire sas_m54;
    reg [63:0] spc54_phy_pc_w;

    

    reg spc55_inst_done;
    wire [1:0]   spc55_thread_id;
    wire [63:0]      spc55_rtl_pc;
    wire sas_m55;
    reg [63:0] spc55_phy_pc_w;

    

    reg spc56_inst_done;
    wire [1:0]   spc56_thread_id;
    wire [63:0]      spc56_rtl_pc;
    wire sas_m56;
    reg [63:0] spc56_phy_pc_w;

    

    reg spc57_inst_done;
    wire [1:0]   spc57_thread_id;
    wire [63:0]      spc57_rtl_pc;
    wire sas_m57;
    reg [63:0] spc57_phy_pc_w;

    

    reg spc58_inst_done;
    wire [1:0]   spc58_thread_id;
    wire [63:0]      spc58_rtl_pc;
    wire sas_m58;
    reg [63:0] spc58_phy_pc_w;

    

    reg spc59_inst_done;
    wire [1:0]   spc59_thread_id;
    wire [63:0]      spc59_rtl_pc;
    wire sas_m59;
    reg [63:0] spc59_phy_pc_w;

    

    reg spc60_inst_done;
    wire [1:0]   spc60_thread_id;
    wire [63:0]      spc60_rtl_pc;
    wire sas_m60;
    reg [63:0] spc60_phy_pc_w;

    

    reg spc61_inst_done;
    wire [1:0]   spc61_thread_id;
    wire [63:0]      spc61_rtl_pc;
    wire sas_m61;
    reg [63:0] spc61_phy_pc_w;

    

    reg spc62_inst_done;
    wire [1:0]   spc62_thread_id;
    wire [63:0]      spc62_rtl_pc;
    wire sas_m62;
    reg [63:0] spc62_phy_pc_w;

    

    reg spc63_inst_done;
    wire [1:0]   spc63_thread_id;
    wire [63:0]      spc63_rtl_pc;
    wire sas_m63;
    reg [63:0] spc63_phy_pc_w;

    

    reg spc64_inst_done;
    wire [1:0]   spc64_thread_id;
    wire [63:0]      spc64_rtl_pc;
    wire sas_m64;
    reg [63:0] spc64_phy_pc_w;

    

    reg spc65_inst_done;
    wire [1:0]   spc65_thread_id;
    wire [63:0]      spc65_rtl_pc;
    wire sas_m65;
    reg [63:0] spc65_phy_pc_w;

    

    reg spc66_inst_done;
    wire [1:0]   spc66_thread_id;
    wire [63:0]      spc66_rtl_pc;
    wire sas_m66;
    reg [63:0] spc66_phy_pc_w;

    

    reg spc67_inst_done;
    wire [1:0]   spc67_thread_id;
    wire [63:0]      spc67_rtl_pc;
    wire sas_m67;
    reg [63:0] spc67_phy_pc_w;

    

    reg spc68_inst_done;
    wire [1:0]   spc68_thread_id;
    wire [63:0]      spc68_rtl_pc;
    wire sas_m68;
    reg [63:0] spc68_phy_pc_w;

    

    reg spc69_inst_done;
    wire [1:0]   spc69_thread_id;
    wire [63:0]      spc69_rtl_pc;
    wire sas_m69;
    reg [63:0] spc69_phy_pc_w;

    

    reg spc70_inst_done;
    wire [1:0]   spc70_thread_id;
    wire [63:0]      spc70_rtl_pc;
    wire sas_m70;
    reg [63:0] spc70_phy_pc_w;

    

    reg spc71_inst_done;
    wire [1:0]   spc71_thread_id;
    wire [63:0]      spc71_rtl_pc;
    wire sas_m71;
    reg [63:0] spc71_phy_pc_w;

    

    reg spc72_inst_done;
    wire [1:0]   spc72_thread_id;
    wire [63:0]      spc72_rtl_pc;
    wire sas_m72;
    reg [63:0] spc72_phy_pc_w;

    

    reg spc73_inst_done;
    wire [1:0]   spc73_thread_id;
    wire [63:0]      spc73_rtl_pc;
    wire sas_m73;
    reg [63:0] spc73_phy_pc_w;

    

    reg spc74_inst_done;
    wire [1:0]   spc74_thread_id;
    wire [63:0]      spc74_rtl_pc;
    wire sas_m74;
    reg [63:0] spc74_phy_pc_w;

    

    reg spc75_inst_done;
    wire [1:0]   spc75_thread_id;
    wire [63:0]      spc75_rtl_pc;
    wire sas_m75;
    reg [63:0] spc75_phy_pc_w;

    

    reg spc76_inst_done;
    wire [1:0]   spc76_thread_id;
    wire [63:0]      spc76_rtl_pc;
    wire sas_m76;
    reg [63:0] spc76_phy_pc_w;

    

    reg spc77_inst_done;
    wire [1:0]   spc77_thread_id;
    wire [63:0]      spc77_rtl_pc;
    wire sas_m77;
    reg [63:0] spc77_phy_pc_w;

    

    reg spc78_inst_done;
    wire [1:0]   spc78_thread_id;
    wire [63:0]      spc78_rtl_pc;
    wire sas_m78;
    reg [63:0] spc78_phy_pc_w;

    

    reg spc79_inst_done;
    wire [1:0]   spc79_thread_id;
    wire [63:0]      spc79_rtl_pc;
    wire sas_m79;
    reg [63:0] spc79_phy_pc_w;

    

    reg spc80_inst_done;
    wire [1:0]   spc80_thread_id;
    wire [63:0]      spc80_rtl_pc;
    wire sas_m80;
    reg [63:0] spc80_phy_pc_w;

    

    reg spc81_inst_done;
    wire [1:0]   spc81_thread_id;
    wire [63:0]      spc81_rtl_pc;
    wire sas_m81;
    reg [63:0] spc81_phy_pc_w;

    

    reg spc82_inst_done;
    wire [1:0]   spc82_thread_id;
    wire [63:0]      spc82_rtl_pc;
    wire sas_m82;
    reg [63:0] spc82_phy_pc_w;

    

    reg spc83_inst_done;
    wire [1:0]   spc83_thread_id;
    wire [63:0]      spc83_rtl_pc;
    wire sas_m83;
    reg [63:0] spc83_phy_pc_w;

    

    reg spc84_inst_done;
    wire [1:0]   spc84_thread_id;
    wire [63:0]      spc84_rtl_pc;
    wire sas_m84;
    reg [63:0] spc84_phy_pc_w;

    

    reg spc85_inst_done;
    wire [1:0]   spc85_thread_id;
    wire [63:0]      spc85_rtl_pc;
    wire sas_m85;
    reg [63:0] spc85_phy_pc_w;

    

    reg spc86_inst_done;
    wire [1:0]   spc86_thread_id;
    wire [63:0]      spc86_rtl_pc;
    wire sas_m86;
    reg [63:0] spc86_phy_pc_w;

    

    reg spc87_inst_done;
    wire [1:0]   spc87_thread_id;
    wire [63:0]      spc87_rtl_pc;
    wire sas_m87;
    reg [63:0] spc87_phy_pc_w;

    

    reg spc88_inst_done;
    wire [1:0]   spc88_thread_id;
    wire [63:0]      spc88_rtl_pc;
    wire sas_m88;
    reg [63:0] spc88_phy_pc_w;

    

    reg spc89_inst_done;
    wire [1:0]   spc89_thread_id;
    wire [63:0]      spc89_rtl_pc;
    wire sas_m89;
    reg [63:0] spc89_phy_pc_w;

    

    reg spc90_inst_done;
    wire [1:0]   spc90_thread_id;
    wire [63:0]      spc90_rtl_pc;
    wire sas_m90;
    reg [63:0] spc90_phy_pc_w;

    

    reg spc91_inst_done;
    wire [1:0]   spc91_thread_id;
    wire [63:0]      spc91_rtl_pc;
    wire sas_m91;
    reg [63:0] spc91_phy_pc_w;

    

    reg spc92_inst_done;
    wire [1:0]   spc92_thread_id;
    wire [63:0]      spc92_rtl_pc;
    wire sas_m92;
    reg [63:0] spc92_phy_pc_w;

    

    reg spc93_inst_done;
    wire [1:0]   spc93_thread_id;
    wire [63:0]      spc93_rtl_pc;
    wire sas_m93;
    reg [63:0] spc93_phy_pc_w;

    

    reg spc94_inst_done;
    wire [1:0]   spc94_thread_id;
    wire [63:0]      spc94_rtl_pc;
    wire sas_m94;
    reg [63:0] spc94_phy_pc_w;

    

    reg spc95_inst_done;
    wire [1:0]   spc95_thread_id;
    wire [63:0]      spc95_rtl_pc;
    wire sas_m95;
    reg [63:0] spc95_phy_pc_w;

    

    reg spc96_inst_done;
    wire [1:0]   spc96_thread_id;
    wire [63:0]      spc96_rtl_pc;
    wire sas_m96;
    reg [63:0] spc96_phy_pc_w;

    

    reg spc97_inst_done;
    wire [1:0]   spc97_thread_id;
    wire [63:0]      spc97_rtl_pc;
    wire sas_m97;
    reg [63:0] spc97_phy_pc_w;

    

    reg spc98_inst_done;
    wire [1:0]   spc98_thread_id;
    wire [63:0]      spc98_rtl_pc;
    wire sas_m98;
    reg [63:0] spc98_phy_pc_w;

    

    reg spc99_inst_done;
    wire [1:0]   spc99_thread_id;
    wire [63:0]      spc99_rtl_pc;
    wire sas_m99;
    reg [63:0] spc99_phy_pc_w;

    

    reg spc100_inst_done;
    wire [1:0]   spc100_thread_id;
    wire [63:0]      spc100_rtl_pc;
    wire sas_m100;
    reg [63:0] spc100_phy_pc_w;

    

    reg spc101_inst_done;
    wire [1:0]   spc101_thread_id;
    wire [63:0]      spc101_rtl_pc;
    wire sas_m101;
    reg [63:0] spc101_phy_pc_w;

    

    reg spc102_inst_done;
    wire [1:0]   spc102_thread_id;
    wire [63:0]      spc102_rtl_pc;
    wire sas_m102;
    reg [63:0] spc102_phy_pc_w;

    

    reg spc103_inst_done;
    wire [1:0]   spc103_thread_id;
    wire [63:0]      spc103_rtl_pc;
    wire sas_m103;
    reg [63:0] spc103_phy_pc_w;

    

    reg spc104_inst_done;
    wire [1:0]   spc104_thread_id;
    wire [63:0]      spc104_rtl_pc;
    wire sas_m104;
    reg [63:0] spc104_phy_pc_w;

    

    reg spc105_inst_done;
    wire [1:0]   spc105_thread_id;
    wire [63:0]      spc105_rtl_pc;
    wire sas_m105;
    reg [63:0] spc105_phy_pc_w;

    

    reg spc106_inst_done;
    wire [1:0]   spc106_thread_id;
    wire [63:0]      spc106_rtl_pc;
    wire sas_m106;
    reg [63:0] spc106_phy_pc_w;

    

    reg spc107_inst_done;
    wire [1:0]   spc107_thread_id;
    wire [63:0]      spc107_rtl_pc;
    wire sas_m107;
    reg [63:0] spc107_phy_pc_w;

    

    reg spc108_inst_done;
    wire [1:0]   spc108_thread_id;
    wire [63:0]      spc108_rtl_pc;
    wire sas_m108;
    reg [63:0] spc108_phy_pc_w;

    

    reg spc109_inst_done;
    wire [1:0]   spc109_thread_id;
    wire [63:0]      spc109_rtl_pc;
    wire sas_m109;
    reg [63:0] spc109_phy_pc_w;

    

    reg spc110_inst_done;
    wire [1:0]   spc110_thread_id;
    wire [63:0]      spc110_rtl_pc;
    wire sas_m110;
    reg [63:0] spc110_phy_pc_w;

    

    reg spc111_inst_done;
    wire [1:0]   spc111_thread_id;
    wire [63:0]      spc111_rtl_pc;
    wire sas_m111;
    reg [63:0] spc111_phy_pc_w;

    

    reg spc112_inst_done;
    wire [1:0]   spc112_thread_id;
    wire [63:0]      spc112_rtl_pc;
    wire sas_m112;
    reg [63:0] spc112_phy_pc_w;

    

    reg spc113_inst_done;
    wire [1:0]   spc113_thread_id;
    wire [63:0]      spc113_rtl_pc;
    wire sas_m113;
    reg [63:0] spc113_phy_pc_w;

    

    reg spc114_inst_done;
    wire [1:0]   spc114_thread_id;
    wire [63:0]      spc114_rtl_pc;
    wire sas_m114;
    reg [63:0] spc114_phy_pc_w;

    

    reg spc115_inst_done;
    wire [1:0]   spc115_thread_id;
    wire [63:0]      spc115_rtl_pc;
    wire sas_m115;
    reg [63:0] spc115_phy_pc_w;

    

    reg spc116_inst_done;
    wire [1:0]   spc116_thread_id;
    wire [63:0]      spc116_rtl_pc;
    wire sas_m116;
    reg [63:0] spc116_phy_pc_w;

    

    reg spc117_inst_done;
    wire [1:0]   spc117_thread_id;
    wire [63:0]      spc117_rtl_pc;
    wire sas_m117;
    reg [63:0] spc117_phy_pc_w;

    

    reg spc118_inst_done;
    wire [1:0]   spc118_thread_id;
    wire [63:0]      spc118_rtl_pc;
    wire sas_m118;
    reg [63:0] spc118_phy_pc_w;

    

    reg spc119_inst_done;
    wire [1:0]   spc119_thread_id;
    wire [63:0]      spc119_rtl_pc;
    wire sas_m119;
    reg [63:0] spc119_phy_pc_w;

    

    reg spc120_inst_done;
    wire [1:0]   spc120_thread_id;
    wire [63:0]      spc120_rtl_pc;
    wire sas_m120;
    reg [63:0] spc120_phy_pc_w;

    

    reg spc121_inst_done;
    wire [1:0]   spc121_thread_id;
    wire [63:0]      spc121_rtl_pc;
    wire sas_m121;
    reg [63:0] spc121_phy_pc_w;

    

    reg spc122_inst_done;
    wire [1:0]   spc122_thread_id;
    wire [63:0]      spc122_rtl_pc;
    wire sas_m122;
    reg [63:0] spc122_phy_pc_w;

    

    reg spc123_inst_done;
    wire [1:0]   spc123_thread_id;
    wire [63:0]      spc123_rtl_pc;
    wire sas_m123;
    reg [63:0] spc123_phy_pc_w;

    

    reg spc124_inst_done;
    wire [1:0]   spc124_thread_id;
    wire [63:0]      spc124_rtl_pc;
    wire sas_m124;
    reg [63:0] spc124_phy_pc_w;

    

    reg spc125_inst_done;
    wire [1:0]   spc125_thread_id;
    wire [63:0]      spc125_rtl_pc;
    wire sas_m125;
    reg [63:0] spc125_phy_pc_w;

    

    reg spc126_inst_done;
    wire [1:0]   spc126_thread_id;
    wire [63:0]      spc126_rtl_pc;
    wire sas_m126;
    reg [63:0] spc126_phy_pc_w;

    

    reg spc127_inst_done;
    wire [1:0]   spc127_thread_id;
    wire [63:0]      spc127_rtl_pc;
    wire sas_m127;
    reg [63:0] spc127_phy_pc_w;

    

    reg spc128_inst_done;
    wire [1:0]   spc128_thread_id;
    wire [63:0]      spc128_rtl_pc;
    wire sas_m128;
    reg [63:0] spc128_phy_pc_w;

    

    reg spc129_inst_done;
    wire [1:0]   spc129_thread_id;
    wire [63:0]      spc129_rtl_pc;
    wire sas_m129;
    reg [63:0] spc129_phy_pc_w;

    

    reg spc130_inst_done;
    wire [1:0]   spc130_thread_id;
    wire [63:0]      spc130_rtl_pc;
    wire sas_m130;
    reg [63:0] spc130_phy_pc_w;

    

    reg spc131_inst_done;
    wire [1:0]   spc131_thread_id;
    wire [63:0]      spc131_rtl_pc;
    wire sas_m131;
    reg [63:0] spc131_phy_pc_w;

    

    reg spc132_inst_done;
    wire [1:0]   spc132_thread_id;
    wire [63:0]      spc132_rtl_pc;
    wire sas_m132;
    reg [63:0] spc132_phy_pc_w;

    

    reg spc133_inst_done;
    wire [1:0]   spc133_thread_id;
    wire [63:0]      spc133_rtl_pc;
    wire sas_m133;
    reg [63:0] spc133_phy_pc_w;

    

    reg spc134_inst_done;
    wire [1:0]   spc134_thread_id;
    wire [63:0]      spc134_rtl_pc;
    wire sas_m134;
    reg [63:0] spc134_phy_pc_w;

    

    reg spc135_inst_done;
    wire [1:0]   spc135_thread_id;
    wire [63:0]      spc135_rtl_pc;
    wire sas_m135;
    reg [63:0] spc135_phy_pc_w;

    

    reg spc136_inst_done;
    wire [1:0]   spc136_thread_id;
    wire [63:0]      spc136_rtl_pc;
    wire sas_m136;
    reg [63:0] spc136_phy_pc_w;

    

    reg spc137_inst_done;
    wire [1:0]   spc137_thread_id;
    wire [63:0]      spc137_rtl_pc;
    wire sas_m137;
    reg [63:0] spc137_phy_pc_w;

    

    reg spc138_inst_done;
    wire [1:0]   spc138_thread_id;
    wire [63:0]      spc138_rtl_pc;
    wire sas_m138;
    reg [63:0] spc138_phy_pc_w;

    

    reg spc139_inst_done;
    wire [1:0]   spc139_thread_id;
    wire [63:0]      spc139_rtl_pc;
    wire sas_m139;
    reg [63:0] spc139_phy_pc_w;

    

    reg spc140_inst_done;
    wire [1:0]   spc140_thread_id;
    wire [63:0]      spc140_rtl_pc;
    wire sas_m140;
    reg [63:0] spc140_phy_pc_w;

    

    reg spc141_inst_done;
    wire [1:0]   spc141_thread_id;
    wire [63:0]      spc141_rtl_pc;
    wire sas_m141;
    reg [63:0] spc141_phy_pc_w;

    

    reg spc142_inst_done;
    wire [1:0]   spc142_thread_id;
    wire [63:0]      spc142_rtl_pc;
    wire sas_m142;
    reg [63:0] spc142_phy_pc_w;

    

    reg spc143_inst_done;
    wire [1:0]   spc143_thread_id;
    wire [63:0]      spc143_rtl_pc;
    wire sas_m143;
    reg [63:0] spc143_phy_pc_w;

    

    reg spc144_inst_done;
    wire [1:0]   spc144_thread_id;
    wire [63:0]      spc144_rtl_pc;
    wire sas_m144;
    reg [63:0] spc144_phy_pc_w;

    

    reg spc145_inst_done;
    wire [1:0]   spc145_thread_id;
    wire [63:0]      spc145_rtl_pc;
    wire sas_m145;
    reg [63:0] spc145_phy_pc_w;

    

    reg spc146_inst_done;
    wire [1:0]   spc146_thread_id;
    wire [63:0]      spc146_rtl_pc;
    wire sas_m146;
    reg [63:0] spc146_phy_pc_w;

    

    reg spc147_inst_done;
    wire [1:0]   spc147_thread_id;
    wire [63:0]      spc147_rtl_pc;
    wire sas_m147;
    reg [63:0] spc147_phy_pc_w;

    

    reg spc148_inst_done;
    wire [1:0]   spc148_thread_id;
    wire [63:0]      spc148_rtl_pc;
    wire sas_m148;
    reg [63:0] spc148_phy_pc_w;

    

    reg spc149_inst_done;
    wire [1:0]   spc149_thread_id;
    wire [63:0]      spc149_rtl_pc;
    wire sas_m149;
    reg [63:0] spc149_phy_pc_w;

    

    reg spc150_inst_done;
    wire [1:0]   spc150_thread_id;
    wire [63:0]      spc150_rtl_pc;
    wire sas_m150;
    reg [63:0] spc150_phy_pc_w;

    

    reg spc151_inst_done;
    wire [1:0]   spc151_thread_id;
    wire [63:0]      spc151_rtl_pc;
    wire sas_m151;
    reg [63:0] spc151_phy_pc_w;

    

    reg spc152_inst_done;
    wire [1:0]   spc152_thread_id;
    wire [63:0]      spc152_rtl_pc;
    wire sas_m152;
    reg [63:0] spc152_phy_pc_w;

    

    reg spc153_inst_done;
    wire [1:0]   spc153_thread_id;
    wire [63:0]      spc153_rtl_pc;
    wire sas_m153;
    reg [63:0] spc153_phy_pc_w;

    

    reg spc154_inst_done;
    wire [1:0]   spc154_thread_id;
    wire [63:0]      spc154_rtl_pc;
    wire sas_m154;
    reg [63:0] spc154_phy_pc_w;

    

    reg spc155_inst_done;
    wire [1:0]   spc155_thread_id;
    wire [63:0]      spc155_rtl_pc;
    wire sas_m155;
    reg [63:0] spc155_phy_pc_w;

    

    reg spc156_inst_done;
    wire [1:0]   spc156_thread_id;
    wire [63:0]      spc156_rtl_pc;
    wire sas_m156;
    reg [63:0] spc156_phy_pc_w;

    

    reg spc157_inst_done;
    wire [1:0]   spc157_thread_id;
    wire [63:0]      spc157_rtl_pc;
    wire sas_m157;
    reg [63:0] spc157_phy_pc_w;

    

    reg spc158_inst_done;
    wire [1:0]   spc158_thread_id;
    wire [63:0]      spc158_rtl_pc;
    wire sas_m158;
    reg [63:0] spc158_phy_pc_w;

    

    reg spc159_inst_done;
    wire [1:0]   spc159_thread_id;
    wire [63:0]      spc159_rtl_pc;
    wire sas_m159;
    reg [63:0] spc159_phy_pc_w;

    

    reg spc160_inst_done;
    wire [1:0]   spc160_thread_id;
    wire [63:0]      spc160_rtl_pc;
    wire sas_m160;
    reg [63:0] spc160_phy_pc_w;

    

    reg spc161_inst_done;
    wire [1:0]   spc161_thread_id;
    wire [63:0]      spc161_rtl_pc;
    wire sas_m161;
    reg [63:0] spc161_phy_pc_w;

    

    reg spc162_inst_done;
    wire [1:0]   spc162_thread_id;
    wire [63:0]      spc162_rtl_pc;
    wire sas_m162;
    reg [63:0] spc162_phy_pc_w;

    

    reg spc163_inst_done;
    wire [1:0]   spc163_thread_id;
    wire [63:0]      spc163_rtl_pc;
    wire sas_m163;
    reg [63:0] spc163_phy_pc_w;

    

    reg spc164_inst_done;
    wire [1:0]   spc164_thread_id;
    wire [63:0]      spc164_rtl_pc;
    wire sas_m164;
    reg [63:0] spc164_phy_pc_w;

    

    reg spc165_inst_done;
    wire [1:0]   spc165_thread_id;
    wire [63:0]      spc165_rtl_pc;
    wire sas_m165;
    reg [63:0] spc165_phy_pc_w;

    

    reg spc166_inst_done;
    wire [1:0]   spc166_thread_id;
    wire [63:0]      spc166_rtl_pc;
    wire sas_m166;
    reg [63:0] spc166_phy_pc_w;

    

    reg spc167_inst_done;
    wire [1:0]   spc167_thread_id;
    wire [63:0]      spc167_rtl_pc;
    wire sas_m167;
    reg [63:0] spc167_phy_pc_w;

    

    reg spc168_inst_done;
    wire [1:0]   spc168_thread_id;
    wire [63:0]      spc168_rtl_pc;
    wire sas_m168;
    reg [63:0] spc168_phy_pc_w;

    

    reg spc169_inst_done;
    wire [1:0]   spc169_thread_id;
    wire [63:0]      spc169_rtl_pc;
    wire sas_m169;
    reg [63:0] spc169_phy_pc_w;

    

    reg spc170_inst_done;
    wire [1:0]   spc170_thread_id;
    wire [63:0]      spc170_rtl_pc;
    wire sas_m170;
    reg [63:0] spc170_phy_pc_w;

    

    reg spc171_inst_done;
    wire [1:0]   spc171_thread_id;
    wire [63:0]      spc171_rtl_pc;
    wire sas_m171;
    reg [63:0] spc171_phy_pc_w;

    

    reg spc172_inst_done;
    wire [1:0]   spc172_thread_id;
    wire [63:0]      spc172_rtl_pc;
    wire sas_m172;
    reg [63:0] spc172_phy_pc_w;

    

    reg spc173_inst_done;
    wire [1:0]   spc173_thread_id;
    wire [63:0]      spc173_rtl_pc;
    wire sas_m173;
    reg [63:0] spc173_phy_pc_w;

    

    reg spc174_inst_done;
    wire [1:0]   spc174_thread_id;
    wire [63:0]      spc174_rtl_pc;
    wire sas_m174;
    reg [63:0] spc174_phy_pc_w;

    

    reg spc175_inst_done;
    wire [1:0]   spc175_thread_id;
    wire [63:0]      spc175_rtl_pc;
    wire sas_m175;
    reg [63:0] spc175_phy_pc_w;

    

    reg spc176_inst_done;
    wire [1:0]   spc176_thread_id;
    wire [63:0]      spc176_rtl_pc;
    wire sas_m176;
    reg [63:0] spc176_phy_pc_w;

    

    reg spc177_inst_done;
    wire [1:0]   spc177_thread_id;
    wire [63:0]      spc177_rtl_pc;
    wire sas_m177;
    reg [63:0] spc177_phy_pc_w;

    

    reg spc178_inst_done;
    wire [1:0]   spc178_thread_id;
    wire [63:0]      spc178_rtl_pc;
    wire sas_m178;
    reg [63:0] spc178_phy_pc_w;

    

    reg spc179_inst_done;
    wire [1:0]   spc179_thread_id;
    wire [63:0]      spc179_rtl_pc;
    wire sas_m179;
    reg [63:0] spc179_phy_pc_w;

    

    reg spc180_inst_done;
    wire [1:0]   spc180_thread_id;
    wire [63:0]      spc180_rtl_pc;
    wire sas_m180;
    reg [63:0] spc180_phy_pc_w;

    

    reg spc181_inst_done;
    wire [1:0]   spc181_thread_id;
    wire [63:0]      spc181_rtl_pc;
    wire sas_m181;
    reg [63:0] spc181_phy_pc_w;

    

    reg spc182_inst_done;
    wire [1:0]   spc182_thread_id;
    wire [63:0]      spc182_rtl_pc;
    wire sas_m182;
    reg [63:0] spc182_phy_pc_w;

    

    reg spc183_inst_done;
    wire [1:0]   spc183_thread_id;
    wire [63:0]      spc183_rtl_pc;
    wire sas_m183;
    reg [63:0] spc183_phy_pc_w;

    

    reg spc184_inst_done;
    wire [1:0]   spc184_thread_id;
    wire [63:0]      spc184_rtl_pc;
    wire sas_m184;
    reg [63:0] spc184_phy_pc_w;

    

    reg spc185_inst_done;
    wire [1:0]   spc185_thread_id;
    wire [63:0]      spc185_rtl_pc;
    wire sas_m185;
    reg [63:0] spc185_phy_pc_w;

    

    reg spc186_inst_done;
    wire [1:0]   spc186_thread_id;
    wire [63:0]      spc186_rtl_pc;
    wire sas_m186;
    reg [63:0] spc186_phy_pc_w;

    

    reg spc187_inst_done;
    wire [1:0]   spc187_thread_id;
    wire [63:0]      spc187_rtl_pc;
    wire sas_m187;
    reg [63:0] spc187_phy_pc_w;

    

    reg spc188_inst_done;
    wire [1:0]   spc188_thread_id;
    wire [63:0]      spc188_rtl_pc;
    wire sas_m188;
    reg [63:0] spc188_phy_pc_w;

    

    reg spc189_inst_done;
    wire [1:0]   spc189_thread_id;
    wire [63:0]      spc189_rtl_pc;
    wire sas_m189;
    reg [63:0] spc189_phy_pc_w;

    

    reg spc190_inst_done;
    wire [1:0]   spc190_thread_id;
    wire [63:0]      spc190_rtl_pc;
    wire sas_m190;
    reg [63:0] spc190_phy_pc_w;

    

    reg spc191_inst_done;
    wire [1:0]   spc191_thread_id;
    wire [63:0]      spc191_rtl_pc;
    wire sas_m191;
    reg [63:0] spc191_phy_pc_w;

    

    reg spc192_inst_done;
    wire [1:0]   spc192_thread_id;
    wire [63:0]      spc192_rtl_pc;
    wire sas_m192;
    reg [63:0] spc192_phy_pc_w;

    

    reg spc193_inst_done;
    wire [1:0]   spc193_thread_id;
    wire [63:0]      spc193_rtl_pc;
    wire sas_m193;
    reg [63:0] spc193_phy_pc_w;

    

    reg spc194_inst_done;
    wire [1:0]   spc194_thread_id;
    wire [63:0]      spc194_rtl_pc;
    wire sas_m194;
    reg [63:0] spc194_phy_pc_w;

    

    reg spc195_inst_done;
    wire [1:0]   spc195_thread_id;
    wire [63:0]      spc195_rtl_pc;
    wire sas_m195;
    reg [63:0] spc195_phy_pc_w;

    

    reg spc196_inst_done;
    wire [1:0]   spc196_thread_id;
    wire [63:0]      spc196_rtl_pc;
    wire sas_m196;
    reg [63:0] spc196_phy_pc_w;

    

    reg spc197_inst_done;
    wire [1:0]   spc197_thread_id;
    wire [63:0]      spc197_rtl_pc;
    wire sas_m197;
    reg [63:0] spc197_phy_pc_w;

    

    reg spc198_inst_done;
    wire [1:0]   spc198_thread_id;
    wire [63:0]      spc198_rtl_pc;
    wire sas_m198;
    reg [63:0] spc198_phy_pc_w;

    

    reg spc199_inst_done;
    wire [1:0]   spc199_thread_id;
    wire [63:0]      spc199_rtl_pc;
    wire sas_m199;
    reg [63:0] spc199_phy_pc_w;

    

    reg spc200_inst_done;
    wire [1:0]   spc200_thread_id;
    wire [63:0]      spc200_rtl_pc;
    wire sas_m200;
    reg [63:0] spc200_phy_pc_w;

    

    reg spc201_inst_done;
    wire [1:0]   spc201_thread_id;
    wire [63:0]      spc201_rtl_pc;
    wire sas_m201;
    reg [63:0] spc201_phy_pc_w;

    

    reg spc202_inst_done;
    wire [1:0]   spc202_thread_id;
    wire [63:0]      spc202_rtl_pc;
    wire sas_m202;
    reg [63:0] spc202_phy_pc_w;

    

    reg spc203_inst_done;
    wire [1:0]   spc203_thread_id;
    wire [63:0]      spc203_rtl_pc;
    wire sas_m203;
    reg [63:0] spc203_phy_pc_w;

    

    reg spc204_inst_done;
    wire [1:0]   spc204_thread_id;
    wire [63:0]      spc204_rtl_pc;
    wire sas_m204;
    reg [63:0] spc204_phy_pc_w;

    

    reg spc205_inst_done;
    wire [1:0]   spc205_thread_id;
    wire [63:0]      spc205_rtl_pc;
    wire sas_m205;
    reg [63:0] spc205_phy_pc_w;

    

    reg spc206_inst_done;
    wire [1:0]   spc206_thread_id;
    wire [63:0]      spc206_rtl_pc;
    wire sas_m206;
    reg [63:0] spc206_phy_pc_w;

    

    reg spc207_inst_done;
    wire [1:0]   spc207_thread_id;
    wire [63:0]      spc207_rtl_pc;
    wire sas_m207;
    reg [63:0] spc207_phy_pc_w;

    

    reg spc208_inst_done;
    wire [1:0]   spc208_thread_id;
    wire [63:0]      spc208_rtl_pc;
    wire sas_m208;
    reg [63:0] spc208_phy_pc_w;

    

    reg spc209_inst_done;
    wire [1:0]   spc209_thread_id;
    wire [63:0]      spc209_rtl_pc;
    wire sas_m209;
    reg [63:0] spc209_phy_pc_w;

    

    reg spc210_inst_done;
    wire [1:0]   spc210_thread_id;
    wire [63:0]      spc210_rtl_pc;
    wire sas_m210;
    reg [63:0] spc210_phy_pc_w;

    

    reg spc211_inst_done;
    wire [1:0]   spc211_thread_id;
    wire [63:0]      spc211_rtl_pc;
    wire sas_m211;
    reg [63:0] spc211_phy_pc_w;

    

    reg spc212_inst_done;
    wire [1:0]   spc212_thread_id;
    wire [63:0]      spc212_rtl_pc;
    wire sas_m212;
    reg [63:0] spc212_phy_pc_w;

    

    reg spc213_inst_done;
    wire [1:0]   spc213_thread_id;
    wire [63:0]      spc213_rtl_pc;
    wire sas_m213;
    reg [63:0] spc213_phy_pc_w;

    

    reg spc214_inst_done;
    wire [1:0]   spc214_thread_id;
    wire [63:0]      spc214_rtl_pc;
    wire sas_m214;
    reg [63:0] spc214_phy_pc_w;

    

    reg spc215_inst_done;
    wire [1:0]   spc215_thread_id;
    wire [63:0]      spc215_rtl_pc;
    wire sas_m215;
    reg [63:0] spc215_phy_pc_w;

    

    reg spc216_inst_done;
    wire [1:0]   spc216_thread_id;
    wire [63:0]      spc216_rtl_pc;
    wire sas_m216;
    reg [63:0] spc216_phy_pc_w;

    

    reg spc217_inst_done;
    wire [1:0]   spc217_thread_id;
    wire [63:0]      spc217_rtl_pc;
    wire sas_m217;
    reg [63:0] spc217_phy_pc_w;

    

    reg spc218_inst_done;
    wire [1:0]   spc218_thread_id;
    wire [63:0]      spc218_rtl_pc;
    wire sas_m218;
    reg [63:0] spc218_phy_pc_w;

    

    reg spc219_inst_done;
    wire [1:0]   spc219_thread_id;
    wire [63:0]      spc219_rtl_pc;
    wire sas_m219;
    reg [63:0] spc219_phy_pc_w;

    

    reg spc220_inst_done;
    wire [1:0]   spc220_thread_id;
    wire [63:0]      spc220_rtl_pc;
    wire sas_m220;
    reg [63:0] spc220_phy_pc_w;

    

    reg spc221_inst_done;
    wire [1:0]   spc221_thread_id;
    wire [63:0]      spc221_rtl_pc;
    wire sas_m221;
    reg [63:0] spc221_phy_pc_w;

    

    reg spc222_inst_done;
    wire [1:0]   spc222_thread_id;
    wire [63:0]      spc222_rtl_pc;
    wire sas_m222;
    reg [63:0] spc222_phy_pc_w;

    

    reg spc223_inst_done;
    wire [1:0]   spc223_thread_id;
    wire [63:0]      spc223_rtl_pc;
    wire sas_m223;
    reg [63:0] spc223_phy_pc_w;

    

    reg spc224_inst_done;
    wire [1:0]   spc224_thread_id;
    wire [63:0]      spc224_rtl_pc;
    wire sas_m224;
    reg [63:0] spc224_phy_pc_w;

    

    reg spc225_inst_done;
    wire [1:0]   spc225_thread_id;
    wire [63:0]      spc225_rtl_pc;
    wire sas_m225;
    reg [63:0] spc225_phy_pc_w;

    

    reg spc226_inst_done;
    wire [1:0]   spc226_thread_id;
    wire [63:0]      spc226_rtl_pc;
    wire sas_m226;
    reg [63:0] spc226_phy_pc_w;

    

    reg spc227_inst_done;
    wire [1:0]   spc227_thread_id;
    wire [63:0]      spc227_rtl_pc;
    wire sas_m227;
    reg [63:0] spc227_phy_pc_w;

    

    reg spc228_inst_done;
    wire [1:0]   spc228_thread_id;
    wire [63:0]      spc228_rtl_pc;
    wire sas_m228;
    reg [63:0] spc228_phy_pc_w;

    

    reg spc229_inst_done;
    wire [1:0]   spc229_thread_id;
    wire [63:0]      spc229_rtl_pc;
    wire sas_m229;
    reg [63:0] spc229_phy_pc_w;

    

    reg spc230_inst_done;
    wire [1:0]   spc230_thread_id;
    wire [63:0]      spc230_rtl_pc;
    wire sas_m230;
    reg [63:0] spc230_phy_pc_w;

    

    reg spc231_inst_done;
    wire [1:0]   spc231_thread_id;
    wire [63:0]      spc231_rtl_pc;
    wire sas_m231;
    reg [63:0] spc231_phy_pc_w;

    

    reg spc232_inst_done;
    wire [1:0]   spc232_thread_id;
    wire [63:0]      spc232_rtl_pc;
    wire sas_m232;
    reg [63:0] spc232_phy_pc_w;

    

    reg spc233_inst_done;
    wire [1:0]   spc233_thread_id;
    wire [63:0]      spc233_rtl_pc;
    wire sas_m233;
    reg [63:0] spc233_phy_pc_w;

    

    reg spc234_inst_done;
    wire [1:0]   spc234_thread_id;
    wire [63:0]      spc234_rtl_pc;
    wire sas_m234;
    reg [63:0] spc234_phy_pc_w;

    

    reg spc235_inst_done;
    wire [1:0]   spc235_thread_id;
    wire [63:0]      spc235_rtl_pc;
    wire sas_m235;
    reg [63:0] spc235_phy_pc_w;

    

    reg spc236_inst_done;
    wire [1:0]   spc236_thread_id;
    wire [63:0]      spc236_rtl_pc;
    wire sas_m236;
    reg [63:0] spc236_phy_pc_w;

    

    reg spc237_inst_done;
    wire [1:0]   spc237_thread_id;
    wire [63:0]      spc237_rtl_pc;
    wire sas_m237;
    reg [63:0] spc237_phy_pc_w;

    

    reg spc238_inst_done;
    wire [1:0]   spc238_thread_id;
    wire [63:0]      spc238_rtl_pc;
    wire sas_m238;
    reg [63:0] spc238_phy_pc_w;

    

    reg spc239_inst_done;
    wire [1:0]   spc239_thread_id;
    wire [63:0]      spc239_rtl_pc;
    wire sas_m239;
    reg [63:0] spc239_phy_pc_w;

    

    reg spc240_inst_done;
    wire [1:0]   spc240_thread_id;
    wire [63:0]      spc240_rtl_pc;
    wire sas_m240;
    reg [63:0] spc240_phy_pc_w;

    

    reg spc241_inst_done;
    wire [1:0]   spc241_thread_id;
    wire [63:0]      spc241_rtl_pc;
    wire sas_m241;
    reg [63:0] spc241_phy_pc_w;

    

    reg spc242_inst_done;
    wire [1:0]   spc242_thread_id;
    wire [63:0]      spc242_rtl_pc;
    wire sas_m242;
    reg [63:0] spc242_phy_pc_w;

    

    reg spc243_inst_done;
    wire [1:0]   spc243_thread_id;
    wire [63:0]      spc243_rtl_pc;
    wire sas_m243;
    reg [63:0] spc243_phy_pc_w;

    

    reg spc244_inst_done;
    wire [1:0]   spc244_thread_id;
    wire [63:0]      spc244_rtl_pc;
    wire sas_m244;
    reg [63:0] spc244_phy_pc_w;

    

    reg spc245_inst_done;
    wire [1:0]   spc245_thread_id;
    wire [63:0]      spc245_rtl_pc;
    wire sas_m245;
    reg [63:0] spc245_phy_pc_w;

    

    reg spc246_inst_done;
    wire [1:0]   spc246_thread_id;
    wire [63:0]      spc246_rtl_pc;
    wire sas_m246;
    reg [63:0] spc246_phy_pc_w;

    

    reg spc247_inst_done;
    wire [1:0]   spc247_thread_id;
    wire [63:0]      spc247_rtl_pc;
    wire sas_m247;
    reg [63:0] spc247_phy_pc_w;

    

    reg spc248_inst_done;
    wire [1:0]   spc248_thread_id;
    wire [63:0]      spc248_rtl_pc;
    wire sas_m248;
    reg [63:0] spc248_phy_pc_w;

    

    reg spc249_inst_done;
    wire [1:0]   spc249_thread_id;
    wire [63:0]      spc249_rtl_pc;
    wire sas_m249;
    reg [63:0] spc249_phy_pc_w;

    

    reg spc250_inst_done;
    wire [1:0]   spc250_thread_id;
    wire [63:0]      spc250_rtl_pc;
    wire sas_m250;
    reg [63:0] spc250_phy_pc_w;

    

    reg spc251_inst_done;
    wire [1:0]   spc251_thread_id;
    wire [63:0]      spc251_rtl_pc;
    wire sas_m251;
    reg [63:0] spc251_phy_pc_w;

    

    reg spc252_inst_done;
    wire [1:0]   spc252_thread_id;
    wire [63:0]      spc252_rtl_pc;
    wire sas_m252;
    reg [63:0] spc252_phy_pc_w;

    

    reg spc253_inst_done;
    wire [1:0]   spc253_thread_id;
    wire [63:0]      spc253_rtl_pc;
    wire sas_m253;
    reg [63:0] spc253_phy_pc_w;

    

    reg spc254_inst_done;
    wire [1:0]   spc254_thread_id;
    wire [63:0]      spc254_rtl_pc;
    wire sas_m254;
    reg [63:0] spc254_phy_pc_w;

    

    reg spc255_inst_done;
    wire [1:0]   spc255_thread_id;
    wire [63:0]      spc255_rtl_pc;
    wire sas_m255;
    reg [63:0] spc255_phy_pc_w;

    

    reg spc256_inst_done;
    wire [1:0]   spc256_thread_id;
    wire [63:0]      spc256_rtl_pc;
    wire sas_m256;
    reg [63:0] spc256_phy_pc_w;

    

    reg spc257_inst_done;
    wire [1:0]   spc257_thread_id;
    wire [63:0]      spc257_rtl_pc;
    wire sas_m257;
    reg [63:0] spc257_phy_pc_w;

    

    reg spc258_inst_done;
    wire [1:0]   spc258_thread_id;
    wire [63:0]      spc258_rtl_pc;
    wire sas_m258;
    reg [63:0] spc258_phy_pc_w;

    

    reg spc259_inst_done;
    wire [1:0]   spc259_thread_id;
    wire [63:0]      spc259_rtl_pc;
    wire sas_m259;
    reg [63:0] spc259_phy_pc_w;

    

    reg spc260_inst_done;
    wire [1:0]   spc260_thread_id;
    wire [63:0]      spc260_rtl_pc;
    wire sas_m260;
    reg [63:0] spc260_phy_pc_w;

    

    reg spc261_inst_done;
    wire [1:0]   spc261_thread_id;
    wire [63:0]      spc261_rtl_pc;
    wire sas_m261;
    reg [63:0] spc261_phy_pc_w;

    

    reg spc262_inst_done;
    wire [1:0]   spc262_thread_id;
    wire [63:0]      spc262_rtl_pc;
    wire sas_m262;
    reg [63:0] spc262_phy_pc_w;

    

    reg spc263_inst_done;
    wire [1:0]   spc263_thread_id;
    wire [63:0]      spc263_rtl_pc;
    wire sas_m263;
    reg [63:0] spc263_phy_pc_w;

    

    reg spc264_inst_done;
    wire [1:0]   spc264_thread_id;
    wire [63:0]      spc264_rtl_pc;
    wire sas_m264;
    reg [63:0] spc264_phy_pc_w;

    

    reg spc265_inst_done;
    wire [1:0]   spc265_thread_id;
    wire [63:0]      spc265_rtl_pc;
    wire sas_m265;
    reg [63:0] spc265_phy_pc_w;

    

    reg spc266_inst_done;
    wire [1:0]   spc266_thread_id;
    wire [63:0]      spc266_rtl_pc;
    wire sas_m266;
    reg [63:0] spc266_phy_pc_w;

    

    reg spc267_inst_done;
    wire [1:0]   spc267_thread_id;
    wire [63:0]      spc267_rtl_pc;
    wire sas_m267;
    reg [63:0] spc267_phy_pc_w;

    

    reg spc268_inst_done;
    wire [1:0]   spc268_thread_id;
    wire [63:0]      spc268_rtl_pc;
    wire sas_m268;
    reg [63:0] spc268_phy_pc_w;

    

    reg spc269_inst_done;
    wire [1:0]   spc269_thread_id;
    wire [63:0]      spc269_rtl_pc;
    wire sas_m269;
    reg [63:0] spc269_phy_pc_w;

    

    reg spc270_inst_done;
    wire [1:0]   spc270_thread_id;
    wire [63:0]      spc270_rtl_pc;
    wire sas_m270;
    reg [63:0] spc270_phy_pc_w;

    

    reg spc271_inst_done;
    wire [1:0]   spc271_thread_id;
    wire [63:0]      spc271_rtl_pc;
    wire sas_m271;
    reg [63:0] spc271_phy_pc_w;

    

    reg spc272_inst_done;
    wire [1:0]   spc272_thread_id;
    wire [63:0]      spc272_rtl_pc;
    wire sas_m272;
    reg [63:0] spc272_phy_pc_w;

    

    reg spc273_inst_done;
    wire [1:0]   spc273_thread_id;
    wire [63:0]      spc273_rtl_pc;
    wire sas_m273;
    reg [63:0] spc273_phy_pc_w;

    

    reg spc274_inst_done;
    wire [1:0]   spc274_thread_id;
    wire [63:0]      spc274_rtl_pc;
    wire sas_m274;
    reg [63:0] spc274_phy_pc_w;

    

    reg spc275_inst_done;
    wire [1:0]   spc275_thread_id;
    wire [63:0]      spc275_rtl_pc;
    wire sas_m275;
    reg [63:0] spc275_phy_pc_w;

    

    reg spc276_inst_done;
    wire [1:0]   spc276_thread_id;
    wire [63:0]      spc276_rtl_pc;
    wire sas_m276;
    reg [63:0] spc276_phy_pc_w;

    

    reg spc277_inst_done;
    wire [1:0]   spc277_thread_id;
    wire [63:0]      spc277_rtl_pc;
    wire sas_m277;
    reg [63:0] spc277_phy_pc_w;

    

    reg spc278_inst_done;
    wire [1:0]   spc278_thread_id;
    wire [63:0]      spc278_rtl_pc;
    wire sas_m278;
    reg [63:0] spc278_phy_pc_w;

    

    reg spc279_inst_done;
    wire [1:0]   spc279_thread_id;
    wire [63:0]      spc279_rtl_pc;
    wire sas_m279;
    reg [63:0] spc279_phy_pc_w;

    

    reg spc280_inst_done;
    wire [1:0]   spc280_thread_id;
    wire [63:0]      spc280_rtl_pc;
    wire sas_m280;
    reg [63:0] spc280_phy_pc_w;

    

    reg spc281_inst_done;
    wire [1:0]   spc281_thread_id;
    wire [63:0]      spc281_rtl_pc;
    wire sas_m281;
    reg [63:0] spc281_phy_pc_w;

    

    reg spc282_inst_done;
    wire [1:0]   spc282_thread_id;
    wire [63:0]      spc282_rtl_pc;
    wire sas_m282;
    reg [63:0] spc282_phy_pc_w;

    

    reg spc283_inst_done;
    wire [1:0]   spc283_thread_id;
    wire [63:0]      spc283_rtl_pc;
    wire sas_m283;
    reg [63:0] spc283_phy_pc_w;

    

    reg spc284_inst_done;
    wire [1:0]   spc284_thread_id;
    wire [63:0]      spc284_rtl_pc;
    wire sas_m284;
    reg [63:0] spc284_phy_pc_w;

    

    reg spc285_inst_done;
    wire [1:0]   spc285_thread_id;
    wire [63:0]      spc285_rtl_pc;
    wire sas_m285;
    reg [63:0] spc285_phy_pc_w;

    

    reg spc286_inst_done;
    wire [1:0]   spc286_thread_id;
    wire [63:0]      spc286_rtl_pc;
    wire sas_m286;
    reg [63:0] spc286_phy_pc_w;

    

    reg spc287_inst_done;
    wire [1:0]   spc287_thread_id;
    wire [63:0]      spc287_rtl_pc;
    wire sas_m287;
    reg [63:0] spc287_phy_pc_w;

    

    reg spc288_inst_done;
    wire [1:0]   spc288_thread_id;
    wire [63:0]      spc288_rtl_pc;
    wire sas_m288;
    reg [63:0] spc288_phy_pc_w;

    

    reg spc289_inst_done;
    wire [1:0]   spc289_thread_id;
    wire [63:0]      spc289_rtl_pc;
    wire sas_m289;
    reg [63:0] spc289_phy_pc_w;

    

    reg spc290_inst_done;
    wire [1:0]   spc290_thread_id;
    wire [63:0]      spc290_rtl_pc;
    wire sas_m290;
    reg [63:0] spc290_phy_pc_w;

    

    reg spc291_inst_done;
    wire [1:0]   spc291_thread_id;
    wire [63:0]      spc291_rtl_pc;
    wire sas_m291;
    reg [63:0] spc291_phy_pc_w;

    

    reg spc292_inst_done;
    wire [1:0]   spc292_thread_id;
    wire [63:0]      spc292_rtl_pc;
    wire sas_m292;
    reg [63:0] spc292_phy_pc_w;

    

    reg spc293_inst_done;
    wire [1:0]   spc293_thread_id;
    wire [63:0]      spc293_rtl_pc;
    wire sas_m293;
    reg [63:0] spc293_phy_pc_w;

    

    reg spc294_inst_done;
    wire [1:0]   spc294_thread_id;
    wire [63:0]      spc294_rtl_pc;
    wire sas_m294;
    reg [63:0] spc294_phy_pc_w;

    

    reg spc295_inst_done;
    wire [1:0]   spc295_thread_id;
    wire [63:0]      spc295_rtl_pc;
    wire sas_m295;
    reg [63:0] spc295_phy_pc_w;

    

    reg spc296_inst_done;
    wire [1:0]   spc296_thread_id;
    wire [63:0]      spc296_rtl_pc;
    wire sas_m296;
    reg [63:0] spc296_phy_pc_w;

    

    reg spc297_inst_done;
    wire [1:0]   spc297_thread_id;
    wire [63:0]      spc297_rtl_pc;
    wire sas_m297;
    reg [63:0] spc297_phy_pc_w;

    

    reg spc298_inst_done;
    wire [1:0]   spc298_thread_id;
    wire [63:0]      spc298_rtl_pc;
    wire sas_m298;
    reg [63:0] spc298_phy_pc_w;

    

    reg spc299_inst_done;
    wire [1:0]   spc299_thread_id;
    wire [63:0]      spc299_rtl_pc;
    wire sas_m299;
    reg [63:0] spc299_phy_pc_w;

    

    reg spc300_inst_done;
    wire [1:0]   spc300_thread_id;
    wire [63:0]      spc300_rtl_pc;
    wire sas_m300;
    reg [63:0] spc300_phy_pc_w;

    

    reg spc301_inst_done;
    wire [1:0]   spc301_thread_id;
    wire [63:0]      spc301_rtl_pc;
    wire sas_m301;
    reg [63:0] spc301_phy_pc_w;

    

    reg spc302_inst_done;
    wire [1:0]   spc302_thread_id;
    wire [63:0]      spc302_rtl_pc;
    wire sas_m302;
    reg [63:0] spc302_phy_pc_w;

    

    reg spc303_inst_done;
    wire [1:0]   spc303_thread_id;
    wire [63:0]      spc303_rtl_pc;
    wire sas_m303;
    reg [63:0] spc303_phy_pc_w;

    

    reg spc304_inst_done;
    wire [1:0]   spc304_thread_id;
    wire [63:0]      spc304_rtl_pc;
    wire sas_m304;
    reg [63:0] spc304_phy_pc_w;

    

    reg spc305_inst_done;
    wire [1:0]   spc305_thread_id;
    wire [63:0]      spc305_rtl_pc;
    wire sas_m305;
    reg [63:0] spc305_phy_pc_w;

    

    reg spc306_inst_done;
    wire [1:0]   spc306_thread_id;
    wire [63:0]      spc306_rtl_pc;
    wire sas_m306;
    reg [63:0] spc306_phy_pc_w;

    

    reg spc307_inst_done;
    wire [1:0]   spc307_thread_id;
    wire [63:0]      spc307_rtl_pc;
    wire sas_m307;
    reg [63:0] spc307_phy_pc_w;

    

    reg spc308_inst_done;
    wire [1:0]   spc308_thread_id;
    wire [63:0]      spc308_rtl_pc;
    wire sas_m308;
    reg [63:0] spc308_phy_pc_w;

    

    reg spc309_inst_done;
    wire [1:0]   spc309_thread_id;
    wire [63:0]      spc309_rtl_pc;
    wire sas_m309;
    reg [63:0] spc309_phy_pc_w;

    

    reg spc310_inst_done;
    wire [1:0]   spc310_thread_id;
    wire [63:0]      spc310_rtl_pc;
    wire sas_m310;
    reg [63:0] spc310_phy_pc_w;

    

    reg spc311_inst_done;
    wire [1:0]   spc311_thread_id;
    wire [63:0]      spc311_rtl_pc;
    wire sas_m311;
    reg [63:0] spc311_phy_pc_w;

    

    reg spc312_inst_done;
    wire [1:0]   spc312_thread_id;
    wire [63:0]      spc312_rtl_pc;
    wire sas_m312;
    reg [63:0] spc312_phy_pc_w;

    

    reg spc313_inst_done;
    wire [1:0]   spc313_thread_id;
    wire [63:0]      spc313_rtl_pc;
    wire sas_m313;
    reg [63:0] spc313_phy_pc_w;

    

    reg spc314_inst_done;
    wire [1:0]   spc314_thread_id;
    wire [63:0]      spc314_rtl_pc;
    wire sas_m314;
    reg [63:0] spc314_phy_pc_w;

    

    reg spc315_inst_done;
    wire [1:0]   spc315_thread_id;
    wire [63:0]      spc315_rtl_pc;
    wire sas_m315;
    reg [63:0] spc315_phy_pc_w;

    

    reg spc316_inst_done;
    wire [1:0]   spc316_thread_id;
    wire [63:0]      spc316_rtl_pc;
    wire sas_m316;
    reg [63:0] spc316_phy_pc_w;

    

    reg spc317_inst_done;
    wire [1:0]   spc317_thread_id;
    wire [63:0]      spc317_rtl_pc;
    wire sas_m317;
    reg [63:0] spc317_phy_pc_w;

    

    reg spc318_inst_done;
    wire [1:0]   spc318_thread_id;
    wire [63:0]      spc318_rtl_pc;
    wire sas_m318;
    reg [63:0] spc318_phy_pc_w;

    

    reg spc319_inst_done;
    wire [1:0]   spc319_thread_id;
    wire [63:0]      spc319_rtl_pc;
    wire sas_m319;
    reg [63:0] spc319_phy_pc_w;

    

    reg spc320_inst_done;
    wire [1:0]   spc320_thread_id;
    wire [63:0]      spc320_rtl_pc;
    wire sas_m320;
    reg [63:0] spc320_phy_pc_w;

    

    reg spc321_inst_done;
    wire [1:0]   spc321_thread_id;
    wire [63:0]      spc321_rtl_pc;
    wire sas_m321;
    reg [63:0] spc321_phy_pc_w;

    

    reg spc322_inst_done;
    wire [1:0]   spc322_thread_id;
    wire [63:0]      spc322_rtl_pc;
    wire sas_m322;
    reg [63:0] spc322_phy_pc_w;

    

    reg spc323_inst_done;
    wire [1:0]   spc323_thread_id;
    wire [63:0]      spc323_rtl_pc;
    wire sas_m323;
    reg [63:0] spc323_phy_pc_w;

    

    reg spc324_inst_done;
    wire [1:0]   spc324_thread_id;
    wire [63:0]      spc324_rtl_pc;
    wire sas_m324;
    reg [63:0] spc324_phy_pc_w;

    

    reg spc325_inst_done;
    wire [1:0]   spc325_thread_id;
    wire [63:0]      spc325_rtl_pc;
    wire sas_m325;
    reg [63:0] spc325_phy_pc_w;

    

    reg spc326_inst_done;
    wire [1:0]   spc326_thread_id;
    wire [63:0]      spc326_rtl_pc;
    wire sas_m326;
    reg [63:0] spc326_phy_pc_w;

    

    reg spc327_inst_done;
    wire [1:0]   spc327_thread_id;
    wire [63:0]      spc327_rtl_pc;
    wire sas_m327;
    reg [63:0] spc327_phy_pc_w;

    

    reg spc328_inst_done;
    wire [1:0]   spc328_thread_id;
    wire [63:0]      spc328_rtl_pc;
    wire sas_m328;
    reg [63:0] spc328_phy_pc_w;

    

    reg spc329_inst_done;
    wire [1:0]   spc329_thread_id;
    wire [63:0]      spc329_rtl_pc;
    wire sas_m329;
    reg [63:0] spc329_phy_pc_w;

    

    reg spc330_inst_done;
    wire [1:0]   spc330_thread_id;
    wire [63:0]      spc330_rtl_pc;
    wire sas_m330;
    reg [63:0] spc330_phy_pc_w;

    

    reg spc331_inst_done;
    wire [1:0]   spc331_thread_id;
    wire [63:0]      spc331_rtl_pc;
    wire sas_m331;
    reg [63:0] spc331_phy_pc_w;

    

    reg spc332_inst_done;
    wire [1:0]   spc332_thread_id;
    wire [63:0]      spc332_rtl_pc;
    wire sas_m332;
    reg [63:0] spc332_phy_pc_w;

    

    reg spc333_inst_done;
    wire [1:0]   spc333_thread_id;
    wire [63:0]      spc333_rtl_pc;
    wire sas_m333;
    reg [63:0] spc333_phy_pc_w;

    

    reg spc334_inst_done;
    wire [1:0]   spc334_thread_id;
    wire [63:0]      spc334_rtl_pc;
    wire sas_m334;
    reg [63:0] spc334_phy_pc_w;

    

    reg spc335_inst_done;
    wire [1:0]   spc335_thread_id;
    wire [63:0]      spc335_rtl_pc;
    wire sas_m335;
    reg [63:0] spc335_phy_pc_w;

    

    reg spc336_inst_done;
    wire [1:0]   spc336_thread_id;
    wire [63:0]      spc336_rtl_pc;
    wire sas_m336;
    reg [63:0] spc336_phy_pc_w;

    

    reg spc337_inst_done;
    wire [1:0]   spc337_thread_id;
    wire [63:0]      spc337_rtl_pc;
    wire sas_m337;
    reg [63:0] spc337_phy_pc_w;

    

    reg spc338_inst_done;
    wire [1:0]   spc338_thread_id;
    wire [63:0]      spc338_rtl_pc;
    wire sas_m338;
    reg [63:0] spc338_phy_pc_w;

    

    reg spc339_inst_done;
    wire [1:0]   spc339_thread_id;
    wire [63:0]      spc339_rtl_pc;
    wire sas_m339;
    reg [63:0] spc339_phy_pc_w;

    

    reg spc340_inst_done;
    wire [1:0]   spc340_thread_id;
    wire [63:0]      spc340_rtl_pc;
    wire sas_m340;
    reg [63:0] spc340_phy_pc_w;

    

    reg spc341_inst_done;
    wire [1:0]   spc341_thread_id;
    wire [63:0]      spc341_rtl_pc;
    wire sas_m341;
    reg [63:0] spc341_phy_pc_w;

    

    reg spc342_inst_done;
    wire [1:0]   spc342_thread_id;
    wire [63:0]      spc342_rtl_pc;
    wire sas_m342;
    reg [63:0] spc342_phy_pc_w;

    

    reg spc343_inst_done;
    wire [1:0]   spc343_thread_id;
    wire [63:0]      spc343_rtl_pc;
    wire sas_m343;
    reg [63:0] spc343_phy_pc_w;

    

    reg spc344_inst_done;
    wire [1:0]   spc344_thread_id;
    wire [63:0]      spc344_rtl_pc;
    wire sas_m344;
    reg [63:0] spc344_phy_pc_w;

    

    reg spc345_inst_done;
    wire [1:0]   spc345_thread_id;
    wire [63:0]      spc345_rtl_pc;
    wire sas_m345;
    reg [63:0] spc345_phy_pc_w;

    

    reg spc346_inst_done;
    wire [1:0]   spc346_thread_id;
    wire [63:0]      spc346_rtl_pc;
    wire sas_m346;
    reg [63:0] spc346_phy_pc_w;

    

    reg spc347_inst_done;
    wire [1:0]   spc347_thread_id;
    wire [63:0]      spc347_rtl_pc;
    wire sas_m347;
    reg [63:0] spc347_phy_pc_w;

    

    reg spc348_inst_done;
    wire [1:0]   spc348_thread_id;
    wire [63:0]      spc348_rtl_pc;
    wire sas_m348;
    reg [63:0] spc348_phy_pc_w;

    

    reg spc349_inst_done;
    wire [1:0]   spc349_thread_id;
    wire [63:0]      spc349_rtl_pc;
    wire sas_m349;
    reg [63:0] spc349_phy_pc_w;

    

    reg spc350_inst_done;
    wire [1:0]   spc350_thread_id;
    wire [63:0]      spc350_rtl_pc;
    wire sas_m350;
    reg [63:0] spc350_phy_pc_w;

    

    reg spc351_inst_done;
    wire [1:0]   spc351_thread_id;
    wire [63:0]      spc351_rtl_pc;
    wire sas_m351;
    reg [63:0] spc351_phy_pc_w;

    

    reg spc352_inst_done;
    wire [1:0]   spc352_thread_id;
    wire [63:0]      spc352_rtl_pc;
    wire sas_m352;
    reg [63:0] spc352_phy_pc_w;

    

    reg spc353_inst_done;
    wire [1:0]   spc353_thread_id;
    wire [63:0]      spc353_rtl_pc;
    wire sas_m353;
    reg [63:0] spc353_phy_pc_w;

    

    reg spc354_inst_done;
    wire [1:0]   spc354_thread_id;
    wire [63:0]      spc354_rtl_pc;
    wire sas_m354;
    reg [63:0] spc354_phy_pc_w;

    

    reg spc355_inst_done;
    wire [1:0]   spc355_thread_id;
    wire [63:0]      spc355_rtl_pc;
    wire sas_m355;
    reg [63:0] spc355_phy_pc_w;

    

    reg spc356_inst_done;
    wire [1:0]   spc356_thread_id;
    wire [63:0]      spc356_rtl_pc;
    wire sas_m356;
    reg [63:0] spc356_phy_pc_w;

    

    reg spc357_inst_done;
    wire [1:0]   spc357_thread_id;
    wire [63:0]      spc357_rtl_pc;
    wire sas_m357;
    reg [63:0] spc357_phy_pc_w;

    

    reg spc358_inst_done;
    wire [1:0]   spc358_thread_id;
    wire [63:0]      spc358_rtl_pc;
    wire sas_m358;
    reg [63:0] spc358_phy_pc_w;

    

    reg spc359_inst_done;
    wire [1:0]   spc359_thread_id;
    wire [63:0]      spc359_rtl_pc;
    wire sas_m359;
    reg [63:0] spc359_phy_pc_w;

    

    reg spc360_inst_done;
    wire [1:0]   spc360_thread_id;
    wire [63:0]      spc360_rtl_pc;
    wire sas_m360;
    reg [63:0] spc360_phy_pc_w;

    

    reg spc361_inst_done;
    wire [1:0]   spc361_thread_id;
    wire [63:0]      spc361_rtl_pc;
    wire sas_m361;
    reg [63:0] spc361_phy_pc_w;

    

    reg spc362_inst_done;
    wire [1:0]   spc362_thread_id;
    wire [63:0]      spc362_rtl_pc;
    wire sas_m362;
    reg [63:0] spc362_phy_pc_w;

    

    reg spc363_inst_done;
    wire [1:0]   spc363_thread_id;
    wire [63:0]      spc363_rtl_pc;
    wire sas_m363;
    reg [63:0] spc363_phy_pc_w;

    

    reg spc364_inst_done;
    wire [1:0]   spc364_thread_id;
    wire [63:0]      spc364_rtl_pc;
    wire sas_m364;
    reg [63:0] spc364_phy_pc_w;

    

    reg spc365_inst_done;
    wire [1:0]   spc365_thread_id;
    wire [63:0]      spc365_rtl_pc;
    wire sas_m365;
    reg [63:0] spc365_phy_pc_w;

    

    reg spc366_inst_done;
    wire [1:0]   spc366_thread_id;
    wire [63:0]      spc366_rtl_pc;
    wire sas_m366;
    reg [63:0] spc366_phy_pc_w;

    

    reg spc367_inst_done;
    wire [1:0]   spc367_thread_id;
    wire [63:0]      spc367_rtl_pc;
    wire sas_m367;
    reg [63:0] spc367_phy_pc_w;

    

    reg spc368_inst_done;
    wire [1:0]   spc368_thread_id;
    wire [63:0]      spc368_rtl_pc;
    wire sas_m368;
    reg [63:0] spc368_phy_pc_w;

    

    reg spc369_inst_done;
    wire [1:0]   spc369_thread_id;
    wire [63:0]      spc369_rtl_pc;
    wire sas_m369;
    reg [63:0] spc369_phy_pc_w;

    

    reg spc370_inst_done;
    wire [1:0]   spc370_thread_id;
    wire [63:0]      spc370_rtl_pc;
    wire sas_m370;
    reg [63:0] spc370_phy_pc_w;

    

    reg spc371_inst_done;
    wire [1:0]   spc371_thread_id;
    wire [63:0]      spc371_rtl_pc;
    wire sas_m371;
    reg [63:0] spc371_phy_pc_w;

    

    reg spc372_inst_done;
    wire [1:0]   spc372_thread_id;
    wire [63:0]      spc372_rtl_pc;
    wire sas_m372;
    reg [63:0] spc372_phy_pc_w;

    

    reg spc373_inst_done;
    wire [1:0]   spc373_thread_id;
    wire [63:0]      spc373_rtl_pc;
    wire sas_m373;
    reg [63:0] spc373_phy_pc_w;

    

    reg spc374_inst_done;
    wire [1:0]   spc374_thread_id;
    wire [63:0]      spc374_rtl_pc;
    wire sas_m374;
    reg [63:0] spc374_phy_pc_w;

    

    reg spc375_inst_done;
    wire [1:0]   spc375_thread_id;
    wire [63:0]      spc375_rtl_pc;
    wire sas_m375;
    reg [63:0] spc375_phy_pc_w;

    

    reg spc376_inst_done;
    wire [1:0]   spc376_thread_id;
    wire [63:0]      spc376_rtl_pc;
    wire sas_m376;
    reg [63:0] spc376_phy_pc_w;

    

    reg spc377_inst_done;
    wire [1:0]   spc377_thread_id;
    wire [63:0]      spc377_rtl_pc;
    wire sas_m377;
    reg [63:0] spc377_phy_pc_w;

    

    reg spc378_inst_done;
    wire [1:0]   spc378_thread_id;
    wire [63:0]      spc378_rtl_pc;
    wire sas_m378;
    reg [63:0] spc378_phy_pc_w;

    

    reg spc379_inst_done;
    wire [1:0]   spc379_thread_id;
    wire [63:0]      spc379_rtl_pc;
    wire sas_m379;
    reg [63:0] spc379_phy_pc_w;

    

    reg spc380_inst_done;
    wire [1:0]   spc380_thread_id;
    wire [63:0]      spc380_rtl_pc;
    wire sas_m380;
    reg [63:0] spc380_phy_pc_w;

    

    reg spc381_inst_done;
    wire [1:0]   spc381_thread_id;
    wire [63:0]      spc381_rtl_pc;
    wire sas_m381;
    reg [63:0] spc381_phy_pc_w;

    

    reg spc382_inst_done;
    wire [1:0]   spc382_thread_id;
    wire [63:0]      spc382_rtl_pc;
    wire sas_m382;
    reg [63:0] spc382_phy_pc_w;

    

    reg spc383_inst_done;
    wire [1:0]   spc383_thread_id;
    wire [63:0]      spc383_rtl_pc;
    wire sas_m383;
    reg [63:0] spc383_phy_pc_w;

    

    reg spc384_inst_done;
    wire [1:0]   spc384_thread_id;
    wire [63:0]      spc384_rtl_pc;
    wire sas_m384;
    reg [63:0] spc384_phy_pc_w;

    

    reg spc385_inst_done;
    wire [1:0]   spc385_thread_id;
    wire [63:0]      spc385_rtl_pc;
    wire sas_m385;
    reg [63:0] spc385_phy_pc_w;

    

    reg spc386_inst_done;
    wire [1:0]   spc386_thread_id;
    wire [63:0]      spc386_rtl_pc;
    wire sas_m386;
    reg [63:0] spc386_phy_pc_w;

    

    reg spc387_inst_done;
    wire [1:0]   spc387_thread_id;
    wire [63:0]      spc387_rtl_pc;
    wire sas_m387;
    reg [63:0] spc387_phy_pc_w;

    

    reg spc388_inst_done;
    wire [1:0]   spc388_thread_id;
    wire [63:0]      spc388_rtl_pc;
    wire sas_m388;
    reg [63:0] spc388_phy_pc_w;

    

    reg spc389_inst_done;
    wire [1:0]   spc389_thread_id;
    wire [63:0]      spc389_rtl_pc;
    wire sas_m389;
    reg [63:0] spc389_phy_pc_w;

    

    reg spc390_inst_done;
    wire [1:0]   spc390_thread_id;
    wire [63:0]      spc390_rtl_pc;
    wire sas_m390;
    reg [63:0] spc390_phy_pc_w;

    

    reg spc391_inst_done;
    wire [1:0]   spc391_thread_id;
    wire [63:0]      spc391_rtl_pc;
    wire sas_m391;
    reg [63:0] spc391_phy_pc_w;

    

    reg spc392_inst_done;
    wire [1:0]   spc392_thread_id;
    wire [63:0]      spc392_rtl_pc;
    wire sas_m392;
    reg [63:0] spc392_phy_pc_w;

    

    reg spc393_inst_done;
    wire [1:0]   spc393_thread_id;
    wire [63:0]      spc393_rtl_pc;
    wire sas_m393;
    reg [63:0] spc393_phy_pc_w;

    

    reg spc394_inst_done;
    wire [1:0]   spc394_thread_id;
    wire [63:0]      spc394_rtl_pc;
    wire sas_m394;
    reg [63:0] spc394_phy_pc_w;

    

    reg spc395_inst_done;
    wire [1:0]   spc395_thread_id;
    wire [63:0]      spc395_rtl_pc;
    wire sas_m395;
    reg [63:0] spc395_phy_pc_w;

    

    reg spc396_inst_done;
    wire [1:0]   spc396_thread_id;
    wire [63:0]      spc396_rtl_pc;
    wire sas_m396;
    reg [63:0] spc396_phy_pc_w;

    

    reg spc397_inst_done;
    wire [1:0]   spc397_thread_id;
    wire [63:0]      spc397_rtl_pc;
    wire sas_m397;
    reg [63:0] spc397_phy_pc_w;

    

    reg spc398_inst_done;
    wire [1:0]   spc398_thread_id;
    wire [63:0]      spc398_rtl_pc;
    wire sas_m398;
    reg [63:0] spc398_phy_pc_w;

    

    reg spc399_inst_done;
    wire [1:0]   spc399_thread_id;
    wire [63:0]      spc399_rtl_pc;
    wire sas_m399;
    reg [63:0] spc399_phy_pc_w;

    

    reg spc400_inst_done;
    wire [1:0]   spc400_thread_id;
    wire [63:0]      spc400_rtl_pc;
    wire sas_m400;
    reg [63:0] spc400_phy_pc_w;

    

    reg spc401_inst_done;
    wire [1:0]   spc401_thread_id;
    wire [63:0]      spc401_rtl_pc;
    wire sas_m401;
    reg [63:0] spc401_phy_pc_w;

    

    reg spc402_inst_done;
    wire [1:0]   spc402_thread_id;
    wire [63:0]      spc402_rtl_pc;
    wire sas_m402;
    reg [63:0] spc402_phy_pc_w;

    

    reg spc403_inst_done;
    wire [1:0]   spc403_thread_id;
    wire [63:0]      spc403_rtl_pc;
    wire sas_m403;
    reg [63:0] spc403_phy_pc_w;

    

    reg spc404_inst_done;
    wire [1:0]   spc404_thread_id;
    wire [63:0]      spc404_rtl_pc;
    wire sas_m404;
    reg [63:0] spc404_phy_pc_w;

    

    reg spc405_inst_done;
    wire [1:0]   spc405_thread_id;
    wire [63:0]      spc405_rtl_pc;
    wire sas_m405;
    reg [63:0] spc405_phy_pc_w;

    

    reg spc406_inst_done;
    wire [1:0]   spc406_thread_id;
    wire [63:0]      spc406_rtl_pc;
    wire sas_m406;
    reg [63:0] spc406_phy_pc_w;

    

    reg spc407_inst_done;
    wire [1:0]   spc407_thread_id;
    wire [63:0]      spc407_rtl_pc;
    wire sas_m407;
    reg [63:0] spc407_phy_pc_w;

    

    reg spc408_inst_done;
    wire [1:0]   spc408_thread_id;
    wire [63:0]      spc408_rtl_pc;
    wire sas_m408;
    reg [63:0] spc408_phy_pc_w;

    

    reg spc409_inst_done;
    wire [1:0]   spc409_thread_id;
    wire [63:0]      spc409_rtl_pc;
    wire sas_m409;
    reg [63:0] spc409_phy_pc_w;

    

    reg spc410_inst_done;
    wire [1:0]   spc410_thread_id;
    wire [63:0]      spc410_rtl_pc;
    wire sas_m410;
    reg [63:0] spc410_phy_pc_w;

    

    reg spc411_inst_done;
    wire [1:0]   spc411_thread_id;
    wire [63:0]      spc411_rtl_pc;
    wire sas_m411;
    reg [63:0] spc411_phy_pc_w;

    

    reg spc412_inst_done;
    wire [1:0]   spc412_thread_id;
    wire [63:0]      spc412_rtl_pc;
    wire sas_m412;
    reg [63:0] spc412_phy_pc_w;

    

    reg spc413_inst_done;
    wire [1:0]   spc413_thread_id;
    wire [63:0]      spc413_rtl_pc;
    wire sas_m413;
    reg [63:0] spc413_phy_pc_w;

    

    reg spc414_inst_done;
    wire [1:0]   spc414_thread_id;
    wire [63:0]      spc414_rtl_pc;
    wire sas_m414;
    reg [63:0] spc414_phy_pc_w;

    

    reg spc415_inst_done;
    wire [1:0]   spc415_thread_id;
    wire [63:0]      spc415_rtl_pc;
    wire sas_m415;
    reg [63:0] spc415_phy_pc_w;

    

    reg spc416_inst_done;
    wire [1:0]   spc416_thread_id;
    wire [63:0]      spc416_rtl_pc;
    wire sas_m416;
    reg [63:0] spc416_phy_pc_w;

    

    reg spc417_inst_done;
    wire [1:0]   spc417_thread_id;
    wire [63:0]      spc417_rtl_pc;
    wire sas_m417;
    reg [63:0] spc417_phy_pc_w;

    

    reg spc418_inst_done;
    wire [1:0]   spc418_thread_id;
    wire [63:0]      spc418_rtl_pc;
    wire sas_m418;
    reg [63:0] spc418_phy_pc_w;

    

    reg spc419_inst_done;
    wire [1:0]   spc419_thread_id;
    wire [63:0]      spc419_rtl_pc;
    wire sas_m419;
    reg [63:0] spc419_phy_pc_w;

    

    reg spc420_inst_done;
    wire [1:0]   spc420_thread_id;
    wire [63:0]      spc420_rtl_pc;
    wire sas_m420;
    reg [63:0] spc420_phy_pc_w;

    

    reg spc421_inst_done;
    wire [1:0]   spc421_thread_id;
    wire [63:0]      spc421_rtl_pc;
    wire sas_m421;
    reg [63:0] spc421_phy_pc_w;

    

    reg spc422_inst_done;
    wire [1:0]   spc422_thread_id;
    wire [63:0]      spc422_rtl_pc;
    wire sas_m422;
    reg [63:0] spc422_phy_pc_w;

    

    reg spc423_inst_done;
    wire [1:0]   spc423_thread_id;
    wire [63:0]      spc423_rtl_pc;
    wire sas_m423;
    reg [63:0] spc423_phy_pc_w;

    

    reg spc424_inst_done;
    wire [1:0]   spc424_thread_id;
    wire [63:0]      spc424_rtl_pc;
    wire sas_m424;
    reg [63:0] spc424_phy_pc_w;

    

    reg spc425_inst_done;
    wire [1:0]   spc425_thread_id;
    wire [63:0]      spc425_rtl_pc;
    wire sas_m425;
    reg [63:0] spc425_phy_pc_w;

    

    reg spc426_inst_done;
    wire [1:0]   spc426_thread_id;
    wire [63:0]      spc426_rtl_pc;
    wire sas_m426;
    reg [63:0] spc426_phy_pc_w;

    

    reg spc427_inst_done;
    wire [1:0]   spc427_thread_id;
    wire [63:0]      spc427_rtl_pc;
    wire sas_m427;
    reg [63:0] spc427_phy_pc_w;

    

    reg spc428_inst_done;
    wire [1:0]   spc428_thread_id;
    wire [63:0]      spc428_rtl_pc;
    wire sas_m428;
    reg [63:0] spc428_phy_pc_w;

    

    reg spc429_inst_done;
    wire [1:0]   spc429_thread_id;
    wire [63:0]      spc429_rtl_pc;
    wire sas_m429;
    reg [63:0] spc429_phy_pc_w;

    

    reg spc430_inst_done;
    wire [1:0]   spc430_thread_id;
    wire [63:0]      spc430_rtl_pc;
    wire sas_m430;
    reg [63:0] spc430_phy_pc_w;

    

    reg spc431_inst_done;
    wire [1:0]   spc431_thread_id;
    wire [63:0]      spc431_rtl_pc;
    wire sas_m431;
    reg [63:0] spc431_phy_pc_w;

    

    reg spc432_inst_done;
    wire [1:0]   spc432_thread_id;
    wire [63:0]      spc432_rtl_pc;
    wire sas_m432;
    reg [63:0] spc432_phy_pc_w;

    

    reg spc433_inst_done;
    wire [1:0]   spc433_thread_id;
    wire [63:0]      spc433_rtl_pc;
    wire sas_m433;
    reg [63:0] spc433_phy_pc_w;

    

    reg spc434_inst_done;
    wire [1:0]   spc434_thread_id;
    wire [63:0]      spc434_rtl_pc;
    wire sas_m434;
    reg [63:0] spc434_phy_pc_w;

    

    reg spc435_inst_done;
    wire [1:0]   spc435_thread_id;
    wire [63:0]      spc435_rtl_pc;
    wire sas_m435;
    reg [63:0] spc435_phy_pc_w;

    

    reg spc436_inst_done;
    wire [1:0]   spc436_thread_id;
    wire [63:0]      spc436_rtl_pc;
    wire sas_m436;
    reg [63:0] spc436_phy_pc_w;

    

    reg spc437_inst_done;
    wire [1:0]   spc437_thread_id;
    wire [63:0]      spc437_rtl_pc;
    wire sas_m437;
    reg [63:0] spc437_phy_pc_w;

    

    reg spc438_inst_done;
    wire [1:0]   spc438_thread_id;
    wire [63:0]      spc438_rtl_pc;
    wire sas_m438;
    reg [63:0] spc438_phy_pc_w;

    

    reg spc439_inst_done;
    wire [1:0]   spc439_thread_id;
    wire [63:0]      spc439_rtl_pc;
    wire sas_m439;
    reg [63:0] spc439_phy_pc_w;

    

    reg spc440_inst_done;
    wire [1:0]   spc440_thread_id;
    wire [63:0]      spc440_rtl_pc;
    wire sas_m440;
    reg [63:0] spc440_phy_pc_w;

    

    reg spc441_inst_done;
    wire [1:0]   spc441_thread_id;
    wire [63:0]      spc441_rtl_pc;
    wire sas_m441;
    reg [63:0] spc441_phy_pc_w;

    

    reg spc442_inst_done;
    wire [1:0]   spc442_thread_id;
    wire [63:0]      spc442_rtl_pc;
    wire sas_m442;
    reg [63:0] spc442_phy_pc_w;

    

    reg spc443_inst_done;
    wire [1:0]   spc443_thread_id;
    wire [63:0]      spc443_rtl_pc;
    wire sas_m443;
    reg [63:0] spc443_phy_pc_w;

    

    reg spc444_inst_done;
    wire [1:0]   spc444_thread_id;
    wire [63:0]      spc444_rtl_pc;
    wire sas_m444;
    reg [63:0] spc444_phy_pc_w;

    

    reg spc445_inst_done;
    wire [1:0]   spc445_thread_id;
    wire [63:0]      spc445_rtl_pc;
    wire sas_m445;
    reg [63:0] spc445_phy_pc_w;

    

    reg spc446_inst_done;
    wire [1:0]   spc446_thread_id;
    wire [63:0]      spc446_rtl_pc;
    wire sas_m446;
    reg [63:0] spc446_phy_pc_w;

    

    reg spc447_inst_done;
    wire [1:0]   spc447_thread_id;
    wire [63:0]      spc447_rtl_pc;
    wire sas_m447;
    reg [63:0] spc447_phy_pc_w;

    

    reg spc448_inst_done;
    wire [1:0]   spc448_thread_id;
    wire [63:0]      spc448_rtl_pc;
    wire sas_m448;
    reg [63:0] spc448_phy_pc_w;

    

    reg spc449_inst_done;
    wire [1:0]   spc449_thread_id;
    wire [63:0]      spc449_rtl_pc;
    wire sas_m449;
    reg [63:0] spc449_phy_pc_w;

    

    reg spc450_inst_done;
    wire [1:0]   spc450_thread_id;
    wire [63:0]      spc450_rtl_pc;
    wire sas_m450;
    reg [63:0] spc450_phy_pc_w;

    

    reg spc451_inst_done;
    wire [1:0]   spc451_thread_id;
    wire [63:0]      spc451_rtl_pc;
    wire sas_m451;
    reg [63:0] spc451_phy_pc_w;

    

    reg spc452_inst_done;
    wire [1:0]   spc452_thread_id;
    wire [63:0]      spc452_rtl_pc;
    wire sas_m452;
    reg [63:0] spc452_phy_pc_w;

    

    reg spc453_inst_done;
    wire [1:0]   spc453_thread_id;
    wire [63:0]      spc453_rtl_pc;
    wire sas_m453;
    reg [63:0] spc453_phy_pc_w;

    

    reg spc454_inst_done;
    wire [1:0]   spc454_thread_id;
    wire [63:0]      spc454_rtl_pc;
    wire sas_m454;
    reg [63:0] spc454_phy_pc_w;

    

    reg spc455_inst_done;
    wire [1:0]   spc455_thread_id;
    wire [63:0]      spc455_rtl_pc;
    wire sas_m455;
    reg [63:0] spc455_phy_pc_w;

    

    reg spc456_inst_done;
    wire [1:0]   spc456_thread_id;
    wire [63:0]      spc456_rtl_pc;
    wire sas_m456;
    reg [63:0] spc456_phy_pc_w;

    

    reg spc457_inst_done;
    wire [1:0]   spc457_thread_id;
    wire [63:0]      spc457_rtl_pc;
    wire sas_m457;
    reg [63:0] spc457_phy_pc_w;

    

    reg spc458_inst_done;
    wire [1:0]   spc458_thread_id;
    wire [63:0]      spc458_rtl_pc;
    wire sas_m458;
    reg [63:0] spc458_phy_pc_w;

    

    reg spc459_inst_done;
    wire [1:0]   spc459_thread_id;
    wire [63:0]      spc459_rtl_pc;
    wire sas_m459;
    reg [63:0] spc459_phy_pc_w;

    

    reg spc460_inst_done;
    wire [1:0]   spc460_thread_id;
    wire [63:0]      spc460_rtl_pc;
    wire sas_m460;
    reg [63:0] spc460_phy_pc_w;

    

    reg spc461_inst_done;
    wire [1:0]   spc461_thread_id;
    wire [63:0]      spc461_rtl_pc;
    wire sas_m461;
    reg [63:0] spc461_phy_pc_w;

    

    reg spc462_inst_done;
    wire [1:0]   spc462_thread_id;
    wire [63:0]      spc462_rtl_pc;
    wire sas_m462;
    reg [63:0] spc462_phy_pc_w;

    

    reg spc463_inst_done;
    wire [1:0]   spc463_thread_id;
    wire [63:0]      spc463_rtl_pc;
    wire sas_m463;
    reg [63:0] spc463_phy_pc_w;

    

    reg spc464_inst_done;
    wire [1:0]   spc464_thread_id;
    wire [63:0]      spc464_rtl_pc;
    wire sas_m464;
    reg [63:0] spc464_phy_pc_w;

    

    reg spc465_inst_done;
    wire [1:0]   spc465_thread_id;
    wire [63:0]      spc465_rtl_pc;
    wire sas_m465;
    reg [63:0] spc465_phy_pc_w;

    

    reg spc466_inst_done;
    wire [1:0]   spc466_thread_id;
    wire [63:0]      spc466_rtl_pc;
    wire sas_m466;
    reg [63:0] spc466_phy_pc_w;

    

    reg spc467_inst_done;
    wire [1:0]   spc467_thread_id;
    wire [63:0]      spc467_rtl_pc;
    wire sas_m467;
    reg [63:0] spc467_phy_pc_w;

    

    reg spc468_inst_done;
    wire [1:0]   spc468_thread_id;
    wire [63:0]      spc468_rtl_pc;
    wire sas_m468;
    reg [63:0] spc468_phy_pc_w;

    

    reg spc469_inst_done;
    wire [1:0]   spc469_thread_id;
    wire [63:0]      spc469_rtl_pc;
    wire sas_m469;
    reg [63:0] spc469_phy_pc_w;

    

    reg spc470_inst_done;
    wire [1:0]   spc470_thread_id;
    wire [63:0]      spc470_rtl_pc;
    wire sas_m470;
    reg [63:0] spc470_phy_pc_w;

    

    reg spc471_inst_done;
    wire [1:0]   spc471_thread_id;
    wire [63:0]      spc471_rtl_pc;
    wire sas_m471;
    reg [63:0] spc471_phy_pc_w;

    

    reg spc472_inst_done;
    wire [1:0]   spc472_thread_id;
    wire [63:0]      spc472_rtl_pc;
    wire sas_m472;
    reg [63:0] spc472_phy_pc_w;

    

    reg spc473_inst_done;
    wire [1:0]   spc473_thread_id;
    wire [63:0]      spc473_rtl_pc;
    wire sas_m473;
    reg [63:0] spc473_phy_pc_w;

    

    reg spc474_inst_done;
    wire [1:0]   spc474_thread_id;
    wire [63:0]      spc474_rtl_pc;
    wire sas_m474;
    reg [63:0] spc474_phy_pc_w;

    

    reg spc475_inst_done;
    wire [1:0]   spc475_thread_id;
    wire [63:0]      spc475_rtl_pc;
    wire sas_m475;
    reg [63:0] spc475_phy_pc_w;

    

    reg spc476_inst_done;
    wire [1:0]   spc476_thread_id;
    wire [63:0]      spc476_rtl_pc;
    wire sas_m476;
    reg [63:0] spc476_phy_pc_w;

    

    reg spc477_inst_done;
    wire [1:0]   spc477_thread_id;
    wire [63:0]      spc477_rtl_pc;
    wire sas_m477;
    reg [63:0] spc477_phy_pc_w;

    

    reg spc478_inst_done;
    wire [1:0]   spc478_thread_id;
    wire [63:0]      spc478_rtl_pc;
    wire sas_m478;
    reg [63:0] spc478_phy_pc_w;

    

    reg spc479_inst_done;
    wire [1:0]   spc479_thread_id;
    wire [63:0]      spc479_rtl_pc;
    wire sas_m479;
    reg [63:0] spc479_phy_pc_w;

    

    reg spc480_inst_done;
    wire [1:0]   spc480_thread_id;
    wire [63:0]      spc480_rtl_pc;
    wire sas_m480;
    reg [63:0] spc480_phy_pc_w;

    

    reg spc481_inst_done;
    wire [1:0]   spc481_thread_id;
    wire [63:0]      spc481_rtl_pc;
    wire sas_m481;
    reg [63:0] spc481_phy_pc_w;

    

    reg spc482_inst_done;
    wire [1:0]   spc482_thread_id;
    wire [63:0]      spc482_rtl_pc;
    wire sas_m482;
    reg [63:0] spc482_phy_pc_w;

    

    reg spc483_inst_done;
    wire [1:0]   spc483_thread_id;
    wire [63:0]      spc483_rtl_pc;
    wire sas_m483;
    reg [63:0] spc483_phy_pc_w;

    

    reg spc484_inst_done;
    wire [1:0]   spc484_thread_id;
    wire [63:0]      spc484_rtl_pc;
    wire sas_m484;
    reg [63:0] spc484_phy_pc_w;

    

    reg spc485_inst_done;
    wire [1:0]   spc485_thread_id;
    wire [63:0]      spc485_rtl_pc;
    wire sas_m485;
    reg [63:0] spc485_phy_pc_w;

    

    reg spc486_inst_done;
    wire [1:0]   spc486_thread_id;
    wire [63:0]      spc486_rtl_pc;
    wire sas_m486;
    reg [63:0] spc486_phy_pc_w;

    

    reg spc487_inst_done;
    wire [1:0]   spc487_thread_id;
    wire [63:0]      spc487_rtl_pc;
    wire sas_m487;
    reg [63:0] spc487_phy_pc_w;

    

    reg spc488_inst_done;
    wire [1:0]   spc488_thread_id;
    wire [63:0]      spc488_rtl_pc;
    wire sas_m488;
    reg [63:0] spc488_phy_pc_w;

    

    reg spc489_inst_done;
    wire [1:0]   spc489_thread_id;
    wire [63:0]      spc489_rtl_pc;
    wire sas_m489;
    reg [63:0] spc489_phy_pc_w;

    

    reg spc490_inst_done;
    wire [1:0]   spc490_thread_id;
    wire [63:0]      spc490_rtl_pc;
    wire sas_m490;
    reg [63:0] spc490_phy_pc_w;

    

    reg spc491_inst_done;
    wire [1:0]   spc491_thread_id;
    wire [63:0]      spc491_rtl_pc;
    wire sas_m491;
    reg [63:0] spc491_phy_pc_w;

    

    reg spc492_inst_done;
    wire [1:0]   spc492_thread_id;
    wire [63:0]      spc492_rtl_pc;
    wire sas_m492;
    reg [63:0] spc492_phy_pc_w;

    

    reg spc493_inst_done;
    wire [1:0]   spc493_thread_id;
    wire [63:0]      spc493_rtl_pc;
    wire sas_m493;
    reg [63:0] spc493_phy_pc_w;

    

    reg spc494_inst_done;
    wire [1:0]   spc494_thread_id;
    wire [63:0]      spc494_rtl_pc;
    wire sas_m494;
    reg [63:0] spc494_phy_pc_w;

    

    reg spc495_inst_done;
    wire [1:0]   spc495_thread_id;
    wire [63:0]      spc495_rtl_pc;
    wire sas_m495;
    reg [63:0] spc495_phy_pc_w;

    

    reg spc496_inst_done;
    wire [1:0]   spc496_thread_id;
    wire [63:0]      spc496_rtl_pc;
    wire sas_m496;
    reg [63:0] spc496_phy_pc_w;

    

    reg spc497_inst_done;
    wire [1:0]   spc497_thread_id;
    wire [63:0]      spc497_rtl_pc;
    wire sas_m497;
    reg [63:0] spc497_phy_pc_w;

    

    reg spc498_inst_done;
    wire [1:0]   spc498_thread_id;
    wire [63:0]      spc498_rtl_pc;
    wire sas_m498;
    reg [63:0] spc498_phy_pc_w;

    

    reg spc499_inst_done;
    wire [1:0]   spc499_thread_id;
    wire [63:0]      spc499_rtl_pc;
    wire sas_m499;
    reg [63:0] spc499_phy_pc_w;

    

    reg spc500_inst_done;
    wire [1:0]   spc500_thread_id;
    wire [63:0]      spc500_rtl_pc;
    wire sas_m500;
    reg [63:0] spc500_phy_pc_w;

    

    reg spc501_inst_done;
    wire [1:0]   spc501_thread_id;
    wire [63:0]      spc501_rtl_pc;
    wire sas_m501;
    reg [63:0] spc501_phy_pc_w;

    

    reg spc502_inst_done;
    wire [1:0]   spc502_thread_id;
    wire [63:0]      spc502_rtl_pc;
    wire sas_m502;
    reg [63:0] spc502_phy_pc_w;

    

    reg spc503_inst_done;
    wire [1:0]   spc503_thread_id;
    wire [63:0]      spc503_rtl_pc;
    wire sas_m503;
    reg [63:0] spc503_phy_pc_w;

    

    reg spc504_inst_done;
    wire [1:0]   spc504_thread_id;
    wire [63:0]      spc504_rtl_pc;
    wire sas_m504;
    reg [63:0] spc504_phy_pc_w;

    

    reg spc505_inst_done;
    wire [1:0]   spc505_thread_id;
    wire [63:0]      spc505_rtl_pc;
    wire sas_m505;
    reg [63:0] spc505_phy_pc_w;

    

    reg spc506_inst_done;
    wire [1:0]   spc506_thread_id;
    wire [63:0]      spc506_rtl_pc;
    wire sas_m506;
    reg [63:0] spc506_phy_pc_w;

    

    reg spc507_inst_done;
    wire [1:0]   spc507_thread_id;
    wire [63:0]      spc507_rtl_pc;
    wire sas_m507;
    reg [63:0] spc507_phy_pc_w;

    

    reg spc508_inst_done;
    wire [1:0]   spc508_thread_id;
    wire [63:0]      spc508_rtl_pc;
    wire sas_m508;
    reg [63:0] spc508_phy_pc_w;

    

    reg spc509_inst_done;
    wire [1:0]   spc509_thread_id;
    wire [63:0]      spc509_rtl_pc;
    wire sas_m509;
    reg [63:0] spc509_phy_pc_w;

    

    reg spc510_inst_done;
    wire [1:0]   spc510_thread_id;
    wire [63:0]      spc510_rtl_pc;
    wire sas_m510;
    reg [63:0] spc510_phy_pc_w;

    

    reg spc511_inst_done;
    wire [1:0]   spc511_thread_id;
    wire [63:0]      spc511_rtl_pc;
    wire sas_m511;
    reg [63:0] spc511_phy_pc_w;

    

    reg spc512_inst_done;
    wire [1:0]   spc512_thread_id;
    wire [63:0]      spc512_rtl_pc;
    wire sas_m512;
    reg [63:0] spc512_phy_pc_w;

    

    reg spc513_inst_done;
    wire [1:0]   spc513_thread_id;
    wire [63:0]      spc513_rtl_pc;
    wire sas_m513;
    reg [63:0] spc513_phy_pc_w;

    

    reg spc514_inst_done;
    wire [1:0]   spc514_thread_id;
    wire [63:0]      spc514_rtl_pc;
    wire sas_m514;
    reg [63:0] spc514_phy_pc_w;

    

    reg spc515_inst_done;
    wire [1:0]   spc515_thread_id;
    wire [63:0]      spc515_rtl_pc;
    wire sas_m515;
    reg [63:0] spc515_phy_pc_w;

    

    reg spc516_inst_done;
    wire [1:0]   spc516_thread_id;
    wire [63:0]      spc516_rtl_pc;
    wire sas_m516;
    reg [63:0] spc516_phy_pc_w;

    

    reg spc517_inst_done;
    wire [1:0]   spc517_thread_id;
    wire [63:0]      spc517_rtl_pc;
    wire sas_m517;
    reg [63:0] spc517_phy_pc_w;

    

    reg spc518_inst_done;
    wire [1:0]   spc518_thread_id;
    wire [63:0]      spc518_rtl_pc;
    wire sas_m518;
    reg [63:0] spc518_phy_pc_w;

    

    reg spc519_inst_done;
    wire [1:0]   spc519_thread_id;
    wire [63:0]      spc519_rtl_pc;
    wire sas_m519;
    reg [63:0] spc519_phy_pc_w;

    

    reg spc520_inst_done;
    wire [1:0]   spc520_thread_id;
    wire [63:0]      spc520_rtl_pc;
    wire sas_m520;
    reg [63:0] spc520_phy_pc_w;

    

    reg spc521_inst_done;
    wire [1:0]   spc521_thread_id;
    wire [63:0]      spc521_rtl_pc;
    wire sas_m521;
    reg [63:0] spc521_phy_pc_w;

    

    reg spc522_inst_done;
    wire [1:0]   spc522_thread_id;
    wire [63:0]      spc522_rtl_pc;
    wire sas_m522;
    reg [63:0] spc522_phy_pc_w;

    

    reg spc523_inst_done;
    wire [1:0]   spc523_thread_id;
    wire [63:0]      spc523_rtl_pc;
    wire sas_m523;
    reg [63:0] spc523_phy_pc_w;

    

    reg spc524_inst_done;
    wire [1:0]   spc524_thread_id;
    wire [63:0]      spc524_rtl_pc;
    wire sas_m524;
    reg [63:0] spc524_phy_pc_w;

    

    reg spc525_inst_done;
    wire [1:0]   spc525_thread_id;
    wire [63:0]      spc525_rtl_pc;
    wire sas_m525;
    reg [63:0] spc525_phy_pc_w;

    

    reg spc526_inst_done;
    wire [1:0]   spc526_thread_id;
    wire [63:0]      spc526_rtl_pc;
    wire sas_m526;
    reg [63:0] spc526_phy_pc_w;

    

    reg spc527_inst_done;
    wire [1:0]   spc527_thread_id;
    wire [63:0]      spc527_rtl_pc;
    wire sas_m527;
    reg [63:0] spc527_phy_pc_w;

    

    reg spc528_inst_done;
    wire [1:0]   spc528_thread_id;
    wire [63:0]      spc528_rtl_pc;
    wire sas_m528;
    reg [63:0] spc528_phy_pc_w;

    

    reg spc529_inst_done;
    wire [1:0]   spc529_thread_id;
    wire [63:0]      spc529_rtl_pc;
    wire sas_m529;
    reg [63:0] spc529_phy_pc_w;

    

    reg spc530_inst_done;
    wire [1:0]   spc530_thread_id;
    wire [63:0]      spc530_rtl_pc;
    wire sas_m530;
    reg [63:0] spc530_phy_pc_w;

    

    reg spc531_inst_done;
    wire [1:0]   spc531_thread_id;
    wire [63:0]      spc531_rtl_pc;
    wire sas_m531;
    reg [63:0] spc531_phy_pc_w;

    

    reg spc532_inst_done;
    wire [1:0]   spc532_thread_id;
    wire [63:0]      spc532_rtl_pc;
    wire sas_m532;
    reg [63:0] spc532_phy_pc_w;

    

    reg spc533_inst_done;
    wire [1:0]   spc533_thread_id;
    wire [63:0]      spc533_rtl_pc;
    wire sas_m533;
    reg [63:0] spc533_phy_pc_w;

    

    reg spc534_inst_done;
    wire [1:0]   spc534_thread_id;
    wire [63:0]      spc534_rtl_pc;
    wire sas_m534;
    reg [63:0] spc534_phy_pc_w;

    

    reg spc535_inst_done;
    wire [1:0]   spc535_thread_id;
    wire [63:0]      spc535_rtl_pc;
    wire sas_m535;
    reg [63:0] spc535_phy_pc_w;

    

    reg spc536_inst_done;
    wire [1:0]   spc536_thread_id;
    wire [63:0]      spc536_rtl_pc;
    wire sas_m536;
    reg [63:0] spc536_phy_pc_w;

    

    reg spc537_inst_done;
    wire [1:0]   spc537_thread_id;
    wire [63:0]      spc537_rtl_pc;
    wire sas_m537;
    reg [63:0] spc537_phy_pc_w;

    

    reg spc538_inst_done;
    wire [1:0]   spc538_thread_id;
    wire [63:0]      spc538_rtl_pc;
    wire sas_m538;
    reg [63:0] spc538_phy_pc_w;

    

    reg spc539_inst_done;
    wire [1:0]   spc539_thread_id;
    wire [63:0]      spc539_rtl_pc;
    wire sas_m539;
    reg [63:0] spc539_phy_pc_w;

    

    reg spc540_inst_done;
    wire [1:0]   spc540_thread_id;
    wire [63:0]      spc540_rtl_pc;
    wire sas_m540;
    reg [63:0] spc540_phy_pc_w;

    

    reg spc541_inst_done;
    wire [1:0]   spc541_thread_id;
    wire [63:0]      spc541_rtl_pc;
    wire sas_m541;
    reg [63:0] spc541_phy_pc_w;

    

    reg spc542_inst_done;
    wire [1:0]   spc542_thread_id;
    wire [63:0]      spc542_rtl_pc;
    wire sas_m542;
    reg [63:0] spc542_phy_pc_w;

    

    reg spc543_inst_done;
    wire [1:0]   spc543_thread_id;
    wire [63:0]      spc543_rtl_pc;
    wire sas_m543;
    reg [63:0] spc543_phy_pc_w;

    

    reg spc544_inst_done;
    wire [1:0]   spc544_thread_id;
    wire [63:0]      spc544_rtl_pc;
    wire sas_m544;
    reg [63:0] spc544_phy_pc_w;

    

    reg spc545_inst_done;
    wire [1:0]   spc545_thread_id;
    wire [63:0]      spc545_rtl_pc;
    wire sas_m545;
    reg [63:0] spc545_phy_pc_w;

    

    reg spc546_inst_done;
    wire [1:0]   spc546_thread_id;
    wire [63:0]      spc546_rtl_pc;
    wire sas_m546;
    reg [63:0] spc546_phy_pc_w;

    

    reg spc547_inst_done;
    wire [1:0]   spc547_thread_id;
    wire [63:0]      spc547_rtl_pc;
    wire sas_m547;
    reg [63:0] spc547_phy_pc_w;

    

    reg spc548_inst_done;
    wire [1:0]   spc548_thread_id;
    wire [63:0]      spc548_rtl_pc;
    wire sas_m548;
    reg [63:0] spc548_phy_pc_w;

    

    reg spc549_inst_done;
    wire [1:0]   spc549_thread_id;
    wire [63:0]      spc549_rtl_pc;
    wire sas_m549;
    reg [63:0] spc549_phy_pc_w;

    

    reg spc550_inst_done;
    wire [1:0]   spc550_thread_id;
    wire [63:0]      spc550_rtl_pc;
    wire sas_m550;
    reg [63:0] spc550_phy_pc_w;

    

    reg spc551_inst_done;
    wire [1:0]   spc551_thread_id;
    wire [63:0]      spc551_rtl_pc;
    wire sas_m551;
    reg [63:0] spc551_phy_pc_w;

    

    reg spc552_inst_done;
    wire [1:0]   spc552_thread_id;
    wire [63:0]      spc552_rtl_pc;
    wire sas_m552;
    reg [63:0] spc552_phy_pc_w;

    

    reg spc553_inst_done;
    wire [1:0]   spc553_thread_id;
    wire [63:0]      spc553_rtl_pc;
    wire sas_m553;
    reg [63:0] spc553_phy_pc_w;

    

    reg spc554_inst_done;
    wire [1:0]   spc554_thread_id;
    wire [63:0]      spc554_rtl_pc;
    wire sas_m554;
    reg [63:0] spc554_phy_pc_w;

    

    reg spc555_inst_done;
    wire [1:0]   spc555_thread_id;
    wire [63:0]      spc555_rtl_pc;
    wire sas_m555;
    reg [63:0] spc555_phy_pc_w;

    

    reg spc556_inst_done;
    wire [1:0]   spc556_thread_id;
    wire [63:0]      spc556_rtl_pc;
    wire sas_m556;
    reg [63:0] spc556_phy_pc_w;

    

    reg spc557_inst_done;
    wire [1:0]   spc557_thread_id;
    wire [63:0]      spc557_rtl_pc;
    wire sas_m557;
    reg [63:0] spc557_phy_pc_w;

    

    reg spc558_inst_done;
    wire [1:0]   spc558_thread_id;
    wire [63:0]      spc558_rtl_pc;
    wire sas_m558;
    reg [63:0] spc558_phy_pc_w;

    

    reg spc559_inst_done;
    wire [1:0]   spc559_thread_id;
    wire [63:0]      spc559_rtl_pc;
    wire sas_m559;
    reg [63:0] spc559_phy_pc_w;

    

    reg spc560_inst_done;
    wire [1:0]   spc560_thread_id;
    wire [63:0]      spc560_rtl_pc;
    wire sas_m560;
    reg [63:0] spc560_phy_pc_w;

    

    reg spc561_inst_done;
    wire [1:0]   spc561_thread_id;
    wire [63:0]      spc561_rtl_pc;
    wire sas_m561;
    reg [63:0] spc561_phy_pc_w;

    

    reg spc562_inst_done;
    wire [1:0]   spc562_thread_id;
    wire [63:0]      spc562_rtl_pc;
    wire sas_m562;
    reg [63:0] spc562_phy_pc_w;

    

    reg spc563_inst_done;
    wire [1:0]   spc563_thread_id;
    wire [63:0]      spc563_rtl_pc;
    wire sas_m563;
    reg [63:0] spc563_phy_pc_w;

    

    reg spc564_inst_done;
    wire [1:0]   spc564_thread_id;
    wire [63:0]      spc564_rtl_pc;
    wire sas_m564;
    reg [63:0] spc564_phy_pc_w;

    

    reg spc565_inst_done;
    wire [1:0]   spc565_thread_id;
    wire [63:0]      spc565_rtl_pc;
    wire sas_m565;
    reg [63:0] spc565_phy_pc_w;

    

    reg spc566_inst_done;
    wire [1:0]   spc566_thread_id;
    wire [63:0]      spc566_rtl_pc;
    wire sas_m566;
    reg [63:0] spc566_phy_pc_w;

    

    reg spc567_inst_done;
    wire [1:0]   spc567_thread_id;
    wire [63:0]      spc567_rtl_pc;
    wire sas_m567;
    reg [63:0] spc567_phy_pc_w;

    

    reg spc568_inst_done;
    wire [1:0]   spc568_thread_id;
    wire [63:0]      spc568_rtl_pc;
    wire sas_m568;
    reg [63:0] spc568_phy_pc_w;

    

    reg spc569_inst_done;
    wire [1:0]   spc569_thread_id;
    wire [63:0]      spc569_rtl_pc;
    wire sas_m569;
    reg [63:0] spc569_phy_pc_w;

    

    reg spc570_inst_done;
    wire [1:0]   spc570_thread_id;
    wire [63:0]      spc570_rtl_pc;
    wire sas_m570;
    reg [63:0] spc570_phy_pc_w;

    

    reg spc571_inst_done;
    wire [1:0]   spc571_thread_id;
    wire [63:0]      spc571_rtl_pc;
    wire sas_m571;
    reg [63:0] spc571_phy_pc_w;

    

    reg spc572_inst_done;
    wire [1:0]   spc572_thread_id;
    wire [63:0]      spc572_rtl_pc;
    wire sas_m572;
    reg [63:0] spc572_phy_pc_w;

    

    reg spc573_inst_done;
    wire [1:0]   spc573_thread_id;
    wire [63:0]      spc573_rtl_pc;
    wire sas_m573;
    reg [63:0] spc573_phy_pc_w;

    

    reg spc574_inst_done;
    wire [1:0]   spc574_thread_id;
    wire [63:0]      spc574_rtl_pc;
    wire sas_m574;
    reg [63:0] spc574_phy_pc_w;

    

    reg spc575_inst_done;
    wire [1:0]   spc575_thread_id;
    wire [63:0]      spc575_rtl_pc;
    wire sas_m575;
    reg [63:0] spc575_phy_pc_w;

    

    reg spc576_inst_done;
    wire [1:0]   spc576_thread_id;
    wire [63:0]      spc576_rtl_pc;
    wire sas_m576;
    reg [63:0] spc576_phy_pc_w;

    

    reg spc577_inst_done;
    wire [1:0]   spc577_thread_id;
    wire [63:0]      spc577_rtl_pc;
    wire sas_m577;
    reg [63:0] spc577_phy_pc_w;

    

    reg spc578_inst_done;
    wire [1:0]   spc578_thread_id;
    wire [63:0]      spc578_rtl_pc;
    wire sas_m578;
    reg [63:0] spc578_phy_pc_w;

    

    reg spc579_inst_done;
    wire [1:0]   spc579_thread_id;
    wire [63:0]      spc579_rtl_pc;
    wire sas_m579;
    reg [63:0] spc579_phy_pc_w;

    

    reg spc580_inst_done;
    wire [1:0]   spc580_thread_id;
    wire [63:0]      spc580_rtl_pc;
    wire sas_m580;
    reg [63:0] spc580_phy_pc_w;

    

    reg spc581_inst_done;
    wire [1:0]   spc581_thread_id;
    wire [63:0]      spc581_rtl_pc;
    wire sas_m581;
    reg [63:0] spc581_phy_pc_w;

    

    reg spc582_inst_done;
    wire [1:0]   spc582_thread_id;
    wire [63:0]      spc582_rtl_pc;
    wire sas_m582;
    reg [63:0] spc582_phy_pc_w;

    

    reg spc583_inst_done;
    wire [1:0]   spc583_thread_id;
    wire [63:0]      spc583_rtl_pc;
    wire sas_m583;
    reg [63:0] spc583_phy_pc_w;

    

    reg spc584_inst_done;
    wire [1:0]   spc584_thread_id;
    wire [63:0]      spc584_rtl_pc;
    wire sas_m584;
    reg [63:0] spc584_phy_pc_w;

    

    reg spc585_inst_done;
    wire [1:0]   spc585_thread_id;
    wire [63:0]      spc585_rtl_pc;
    wire sas_m585;
    reg [63:0] spc585_phy_pc_w;

    

    reg spc586_inst_done;
    wire [1:0]   spc586_thread_id;
    wire [63:0]      spc586_rtl_pc;
    wire sas_m586;
    reg [63:0] spc586_phy_pc_w;

    

    reg spc587_inst_done;
    wire [1:0]   spc587_thread_id;
    wire [63:0]      spc587_rtl_pc;
    wire sas_m587;
    reg [63:0] spc587_phy_pc_w;

    

    reg spc588_inst_done;
    wire [1:0]   spc588_thread_id;
    wire [63:0]      spc588_rtl_pc;
    wire sas_m588;
    reg [63:0] spc588_phy_pc_w;

    

    reg spc589_inst_done;
    wire [1:0]   spc589_thread_id;
    wire [63:0]      spc589_rtl_pc;
    wire sas_m589;
    reg [63:0] spc589_phy_pc_w;

    

    reg spc590_inst_done;
    wire [1:0]   spc590_thread_id;
    wire [63:0]      spc590_rtl_pc;
    wire sas_m590;
    reg [63:0] spc590_phy_pc_w;

    

    reg spc591_inst_done;
    wire [1:0]   spc591_thread_id;
    wire [63:0]      spc591_rtl_pc;
    wire sas_m591;
    reg [63:0] spc591_phy_pc_w;

    

    reg spc592_inst_done;
    wire [1:0]   spc592_thread_id;
    wire [63:0]      spc592_rtl_pc;
    wire sas_m592;
    reg [63:0] spc592_phy_pc_w;

    

    reg spc593_inst_done;
    wire [1:0]   spc593_thread_id;
    wire [63:0]      spc593_rtl_pc;
    wire sas_m593;
    reg [63:0] spc593_phy_pc_w;

    

    reg spc594_inst_done;
    wire [1:0]   spc594_thread_id;
    wire [63:0]      spc594_rtl_pc;
    wire sas_m594;
    reg [63:0] spc594_phy_pc_w;

    

    reg spc595_inst_done;
    wire [1:0]   spc595_thread_id;
    wire [63:0]      spc595_rtl_pc;
    wire sas_m595;
    reg [63:0] spc595_phy_pc_w;

    

    reg spc596_inst_done;
    wire [1:0]   spc596_thread_id;
    wire [63:0]      spc596_rtl_pc;
    wire sas_m596;
    reg [63:0] spc596_phy_pc_w;

    

    reg spc597_inst_done;
    wire [1:0]   spc597_thread_id;
    wire [63:0]      spc597_rtl_pc;
    wire sas_m597;
    reg [63:0] spc597_phy_pc_w;

    

    reg spc598_inst_done;
    wire [1:0]   spc598_thread_id;
    wire [63:0]      spc598_rtl_pc;
    wire sas_m598;
    reg [63:0] spc598_phy_pc_w;

    

    reg spc599_inst_done;
    wire [1:0]   spc599_thread_id;
    wire [63:0]      spc599_rtl_pc;
    wire sas_m599;
    reg [63:0] spc599_phy_pc_w;

    

    reg spc600_inst_done;
    wire [1:0]   spc600_thread_id;
    wire [63:0]      spc600_rtl_pc;
    wire sas_m600;
    reg [63:0] spc600_phy_pc_w;

    

    reg spc601_inst_done;
    wire [1:0]   spc601_thread_id;
    wire [63:0]      spc601_rtl_pc;
    wire sas_m601;
    reg [63:0] spc601_phy_pc_w;

    

    reg spc602_inst_done;
    wire [1:0]   spc602_thread_id;
    wire [63:0]      spc602_rtl_pc;
    wire sas_m602;
    reg [63:0] spc602_phy_pc_w;

    

    reg spc603_inst_done;
    wire [1:0]   spc603_thread_id;
    wire [63:0]      spc603_rtl_pc;
    wire sas_m603;
    reg [63:0] spc603_phy_pc_w;

    

    reg spc604_inst_done;
    wire [1:0]   spc604_thread_id;
    wire [63:0]      spc604_rtl_pc;
    wire sas_m604;
    reg [63:0] spc604_phy_pc_w;

    

    reg spc605_inst_done;
    wire [1:0]   spc605_thread_id;
    wire [63:0]      spc605_rtl_pc;
    wire sas_m605;
    reg [63:0] spc605_phy_pc_w;

    

    reg spc606_inst_done;
    wire [1:0]   spc606_thread_id;
    wire [63:0]      spc606_rtl_pc;
    wire sas_m606;
    reg [63:0] spc606_phy_pc_w;

    

    reg spc607_inst_done;
    wire [1:0]   spc607_thread_id;
    wire [63:0]      spc607_rtl_pc;
    wire sas_m607;
    reg [63:0] spc607_phy_pc_w;

    

    reg spc608_inst_done;
    wire [1:0]   spc608_thread_id;
    wire [63:0]      spc608_rtl_pc;
    wire sas_m608;
    reg [63:0] spc608_phy_pc_w;

    

    reg spc609_inst_done;
    wire [1:0]   spc609_thread_id;
    wire [63:0]      spc609_rtl_pc;
    wire sas_m609;
    reg [63:0] spc609_phy_pc_w;

    

    reg spc610_inst_done;
    wire [1:0]   spc610_thread_id;
    wire [63:0]      spc610_rtl_pc;
    wire sas_m610;
    reg [63:0] spc610_phy_pc_w;

    

    reg spc611_inst_done;
    wire [1:0]   spc611_thread_id;
    wire [63:0]      spc611_rtl_pc;
    wire sas_m611;
    reg [63:0] spc611_phy_pc_w;

    

    reg spc612_inst_done;
    wire [1:0]   spc612_thread_id;
    wire [63:0]      spc612_rtl_pc;
    wire sas_m612;
    reg [63:0] spc612_phy_pc_w;

    

    reg spc613_inst_done;
    wire [1:0]   spc613_thread_id;
    wire [63:0]      spc613_rtl_pc;
    wire sas_m613;
    reg [63:0] spc613_phy_pc_w;

    

    reg spc614_inst_done;
    wire [1:0]   spc614_thread_id;
    wire [63:0]      spc614_rtl_pc;
    wire sas_m614;
    reg [63:0] spc614_phy_pc_w;

    

    reg spc615_inst_done;
    wire [1:0]   spc615_thread_id;
    wire [63:0]      spc615_rtl_pc;
    wire sas_m615;
    reg [63:0] spc615_phy_pc_w;

    

    reg spc616_inst_done;
    wire [1:0]   spc616_thread_id;
    wire [63:0]      spc616_rtl_pc;
    wire sas_m616;
    reg [63:0] spc616_phy_pc_w;

    

    reg spc617_inst_done;
    wire [1:0]   spc617_thread_id;
    wire [63:0]      spc617_rtl_pc;
    wire sas_m617;
    reg [63:0] spc617_phy_pc_w;

    

    reg spc618_inst_done;
    wire [1:0]   spc618_thread_id;
    wire [63:0]      spc618_rtl_pc;
    wire sas_m618;
    reg [63:0] spc618_phy_pc_w;

    

    reg spc619_inst_done;
    wire [1:0]   spc619_thread_id;
    wire [63:0]      spc619_rtl_pc;
    wire sas_m619;
    reg [63:0] spc619_phy_pc_w;

    

    reg spc620_inst_done;
    wire [1:0]   spc620_thread_id;
    wire [63:0]      spc620_rtl_pc;
    wire sas_m620;
    reg [63:0] spc620_phy_pc_w;

    

    reg spc621_inst_done;
    wire [1:0]   spc621_thread_id;
    wire [63:0]      spc621_rtl_pc;
    wire sas_m621;
    reg [63:0] spc621_phy_pc_w;

    

    reg spc622_inst_done;
    wire [1:0]   spc622_thread_id;
    wire [63:0]      spc622_rtl_pc;
    wire sas_m622;
    reg [63:0] spc622_phy_pc_w;

    

    reg spc623_inst_done;
    wire [1:0]   spc623_thread_id;
    wire [63:0]      spc623_rtl_pc;
    wire sas_m623;
    reg [63:0] spc623_phy_pc_w;

    

    reg spc624_inst_done;
    wire [1:0]   spc624_thread_id;
    wire [63:0]      spc624_rtl_pc;
    wire sas_m624;
    reg [63:0] spc624_phy_pc_w;

    

    reg spc625_inst_done;
    wire [1:0]   spc625_thread_id;
    wire [63:0]      spc625_rtl_pc;
    wire sas_m625;
    reg [63:0] spc625_phy_pc_w;

    

    reg spc626_inst_done;
    wire [1:0]   spc626_thread_id;
    wire [63:0]      spc626_rtl_pc;
    wire sas_m626;
    reg [63:0] spc626_phy_pc_w;

    

    reg spc627_inst_done;
    wire [1:0]   spc627_thread_id;
    wire [63:0]      spc627_rtl_pc;
    wire sas_m627;
    reg [63:0] spc627_phy_pc_w;

    

    reg spc628_inst_done;
    wire [1:0]   spc628_thread_id;
    wire [63:0]      spc628_rtl_pc;
    wire sas_m628;
    reg [63:0] spc628_phy_pc_w;

    

    reg spc629_inst_done;
    wire [1:0]   spc629_thread_id;
    wire [63:0]      spc629_rtl_pc;
    wire sas_m629;
    reg [63:0] spc629_phy_pc_w;

    

    reg spc630_inst_done;
    wire [1:0]   spc630_thread_id;
    wire [63:0]      spc630_rtl_pc;
    wire sas_m630;
    reg [63:0] spc630_phy_pc_w;

    

    reg spc631_inst_done;
    wire [1:0]   spc631_thread_id;
    wire [63:0]      spc631_rtl_pc;
    wire sas_m631;
    reg [63:0] spc631_phy_pc_w;

    

    reg spc632_inst_done;
    wire [1:0]   spc632_thread_id;
    wire [63:0]      spc632_rtl_pc;
    wire sas_m632;
    reg [63:0] spc632_phy_pc_w;

    

    reg spc633_inst_done;
    wire [1:0]   spc633_thread_id;
    wire [63:0]      spc633_rtl_pc;
    wire sas_m633;
    reg [63:0] spc633_phy_pc_w;

    

    reg spc634_inst_done;
    wire [1:0]   spc634_thread_id;
    wire [63:0]      spc634_rtl_pc;
    wire sas_m634;
    reg [63:0] spc634_phy_pc_w;

    

    reg spc635_inst_done;
    wire [1:0]   spc635_thread_id;
    wire [63:0]      spc635_rtl_pc;
    wire sas_m635;
    reg [63:0] spc635_phy_pc_w;

    

    reg spc636_inst_done;
    wire [1:0]   spc636_thread_id;
    wire [63:0]      spc636_rtl_pc;
    wire sas_m636;
    reg [63:0] spc636_phy_pc_w;

    

    reg spc637_inst_done;
    wire [1:0]   spc637_thread_id;
    wire [63:0]      spc637_rtl_pc;
    wire sas_m637;
    reg [63:0] spc637_phy_pc_w;

    

    reg spc638_inst_done;
    wire [1:0]   spc638_thread_id;
    wire [63:0]      spc638_rtl_pc;
    wire sas_m638;
    reg [63:0] spc638_phy_pc_w;

    

    reg spc639_inst_done;
    wire [1:0]   spc639_thread_id;
    wire [63:0]      spc639_rtl_pc;
    wire sas_m639;
    reg [63:0] spc639_phy_pc_w;

    

    reg spc640_inst_done;
    wire [1:0]   spc640_thread_id;
    wire [63:0]      spc640_rtl_pc;
    wire sas_m640;
    reg [63:0] spc640_phy_pc_w;

    

    reg spc641_inst_done;
    wire [1:0]   spc641_thread_id;
    wire [63:0]      spc641_rtl_pc;
    wire sas_m641;
    reg [63:0] spc641_phy_pc_w;

    

    reg spc642_inst_done;
    wire [1:0]   spc642_thread_id;
    wire [63:0]      spc642_rtl_pc;
    wire sas_m642;
    reg [63:0] spc642_phy_pc_w;

    

    reg spc643_inst_done;
    wire [1:0]   spc643_thread_id;
    wire [63:0]      spc643_rtl_pc;
    wire sas_m643;
    reg [63:0] spc643_phy_pc_w;

    

    reg spc644_inst_done;
    wire [1:0]   spc644_thread_id;
    wire [63:0]      spc644_rtl_pc;
    wire sas_m644;
    reg [63:0] spc644_phy_pc_w;

    

    reg spc645_inst_done;
    wire [1:0]   spc645_thread_id;
    wire [63:0]      spc645_rtl_pc;
    wire sas_m645;
    reg [63:0] spc645_phy_pc_w;

    

    reg spc646_inst_done;
    wire [1:0]   spc646_thread_id;
    wire [63:0]      spc646_rtl_pc;
    wire sas_m646;
    reg [63:0] spc646_phy_pc_w;

    

    reg spc647_inst_done;
    wire [1:0]   spc647_thread_id;
    wire [63:0]      spc647_rtl_pc;
    wire sas_m647;
    reg [63:0] spc647_phy_pc_w;

    

    reg spc648_inst_done;
    wire [1:0]   spc648_thread_id;
    wire [63:0]      spc648_rtl_pc;
    wire sas_m648;
    reg [63:0] spc648_phy_pc_w;

    

    reg spc649_inst_done;
    wire [1:0]   spc649_thread_id;
    wire [63:0]      spc649_rtl_pc;
    wire sas_m649;
    reg [63:0] spc649_phy_pc_w;

    

    reg spc650_inst_done;
    wire [1:0]   spc650_thread_id;
    wire [63:0]      spc650_rtl_pc;
    wire sas_m650;
    reg [63:0] spc650_phy_pc_w;

    

    reg spc651_inst_done;
    wire [1:0]   spc651_thread_id;
    wire [63:0]      spc651_rtl_pc;
    wire sas_m651;
    reg [63:0] spc651_phy_pc_w;

    

    reg spc652_inst_done;
    wire [1:0]   spc652_thread_id;
    wire [63:0]      spc652_rtl_pc;
    wire sas_m652;
    reg [63:0] spc652_phy_pc_w;

    

    reg spc653_inst_done;
    wire [1:0]   spc653_thread_id;
    wire [63:0]      spc653_rtl_pc;
    wire sas_m653;
    reg [63:0] spc653_phy_pc_w;

    

    reg spc654_inst_done;
    wire [1:0]   spc654_thread_id;
    wire [63:0]      spc654_rtl_pc;
    wire sas_m654;
    reg [63:0] spc654_phy_pc_w;

    

    reg spc655_inst_done;
    wire [1:0]   spc655_thread_id;
    wire [63:0]      spc655_rtl_pc;
    wire sas_m655;
    reg [63:0] spc655_phy_pc_w;

    

    reg spc656_inst_done;
    wire [1:0]   spc656_thread_id;
    wire [63:0]      spc656_rtl_pc;
    wire sas_m656;
    reg [63:0] spc656_phy_pc_w;

    

    reg spc657_inst_done;
    wire [1:0]   spc657_thread_id;
    wire [63:0]      spc657_rtl_pc;
    wire sas_m657;
    reg [63:0] spc657_phy_pc_w;

    

    reg spc658_inst_done;
    wire [1:0]   spc658_thread_id;
    wire [63:0]      spc658_rtl_pc;
    wire sas_m658;
    reg [63:0] spc658_phy_pc_w;

    

    reg spc659_inst_done;
    wire [1:0]   spc659_thread_id;
    wire [63:0]      spc659_rtl_pc;
    wire sas_m659;
    reg [63:0] spc659_phy_pc_w;

    

    reg spc660_inst_done;
    wire [1:0]   spc660_thread_id;
    wire [63:0]      spc660_rtl_pc;
    wire sas_m660;
    reg [63:0] spc660_phy_pc_w;

    

    reg spc661_inst_done;
    wire [1:0]   spc661_thread_id;
    wire [63:0]      spc661_rtl_pc;
    wire sas_m661;
    reg [63:0] spc661_phy_pc_w;

    

    reg spc662_inst_done;
    wire [1:0]   spc662_thread_id;
    wire [63:0]      spc662_rtl_pc;
    wire sas_m662;
    reg [63:0] spc662_phy_pc_w;

    

    reg spc663_inst_done;
    wire [1:0]   spc663_thread_id;
    wire [63:0]      spc663_rtl_pc;
    wire sas_m663;
    reg [63:0] spc663_phy_pc_w;

    

    reg spc664_inst_done;
    wire [1:0]   spc664_thread_id;
    wire [63:0]      spc664_rtl_pc;
    wire sas_m664;
    reg [63:0] spc664_phy_pc_w;

    

    reg spc665_inst_done;
    wire [1:0]   spc665_thread_id;
    wire [63:0]      spc665_rtl_pc;
    wire sas_m665;
    reg [63:0] spc665_phy_pc_w;

    

    reg spc666_inst_done;
    wire [1:0]   spc666_thread_id;
    wire [63:0]      spc666_rtl_pc;
    wire sas_m666;
    reg [63:0] spc666_phy_pc_w;

    

    reg spc667_inst_done;
    wire [1:0]   spc667_thread_id;
    wire [63:0]      spc667_rtl_pc;
    wire sas_m667;
    reg [63:0] spc667_phy_pc_w;

    

    reg spc668_inst_done;
    wire [1:0]   spc668_thread_id;
    wire [63:0]      spc668_rtl_pc;
    wire sas_m668;
    reg [63:0] spc668_phy_pc_w;

    

    reg spc669_inst_done;
    wire [1:0]   spc669_thread_id;
    wire [63:0]      spc669_rtl_pc;
    wire sas_m669;
    reg [63:0] spc669_phy_pc_w;

    

    reg spc670_inst_done;
    wire [1:0]   spc670_thread_id;
    wire [63:0]      spc670_rtl_pc;
    wire sas_m670;
    reg [63:0] spc670_phy_pc_w;

    

    reg spc671_inst_done;
    wire [1:0]   spc671_thread_id;
    wire [63:0]      spc671_rtl_pc;
    wire sas_m671;
    reg [63:0] spc671_phy_pc_w;

    

    reg spc672_inst_done;
    wire [1:0]   spc672_thread_id;
    wire [63:0]      spc672_rtl_pc;
    wire sas_m672;
    reg [63:0] spc672_phy_pc_w;

    

    reg spc673_inst_done;
    wire [1:0]   spc673_thread_id;
    wire [63:0]      spc673_rtl_pc;
    wire sas_m673;
    reg [63:0] spc673_phy_pc_w;

    

    reg spc674_inst_done;
    wire [1:0]   spc674_thread_id;
    wire [63:0]      spc674_rtl_pc;
    wire sas_m674;
    reg [63:0] spc674_phy_pc_w;

    

    reg spc675_inst_done;
    wire [1:0]   spc675_thread_id;
    wire [63:0]      spc675_rtl_pc;
    wire sas_m675;
    reg [63:0] spc675_phy_pc_w;

    

    reg spc676_inst_done;
    wire [1:0]   spc676_thread_id;
    wire [63:0]      spc676_rtl_pc;
    wire sas_m676;
    reg [63:0] spc676_phy_pc_w;

    

    reg spc677_inst_done;
    wire [1:0]   spc677_thread_id;
    wire [63:0]      spc677_rtl_pc;
    wire sas_m677;
    reg [63:0] spc677_phy_pc_w;

    

    reg spc678_inst_done;
    wire [1:0]   spc678_thread_id;
    wire [63:0]      spc678_rtl_pc;
    wire sas_m678;
    reg [63:0] spc678_phy_pc_w;

    

    reg spc679_inst_done;
    wire [1:0]   spc679_thread_id;
    wire [63:0]      spc679_rtl_pc;
    wire sas_m679;
    reg [63:0] spc679_phy_pc_w;

    

    reg spc680_inst_done;
    wire [1:0]   spc680_thread_id;
    wire [63:0]      spc680_rtl_pc;
    wire sas_m680;
    reg [63:0] spc680_phy_pc_w;

    

    reg spc681_inst_done;
    wire [1:0]   spc681_thread_id;
    wire [63:0]      spc681_rtl_pc;
    wire sas_m681;
    reg [63:0] spc681_phy_pc_w;

    

    reg spc682_inst_done;
    wire [1:0]   spc682_thread_id;
    wire [63:0]      spc682_rtl_pc;
    wire sas_m682;
    reg [63:0] spc682_phy_pc_w;

    

    reg spc683_inst_done;
    wire [1:0]   spc683_thread_id;
    wire [63:0]      spc683_rtl_pc;
    wire sas_m683;
    reg [63:0] spc683_phy_pc_w;

    

    reg spc684_inst_done;
    wire [1:0]   spc684_thread_id;
    wire [63:0]      spc684_rtl_pc;
    wire sas_m684;
    reg [63:0] spc684_phy_pc_w;

    

    reg spc685_inst_done;
    wire [1:0]   spc685_thread_id;
    wire [63:0]      spc685_rtl_pc;
    wire sas_m685;
    reg [63:0] spc685_phy_pc_w;

    

    reg spc686_inst_done;
    wire [1:0]   spc686_thread_id;
    wire [63:0]      spc686_rtl_pc;
    wire sas_m686;
    reg [63:0] spc686_phy_pc_w;

    

    reg spc687_inst_done;
    wire [1:0]   spc687_thread_id;
    wire [63:0]      spc687_rtl_pc;
    wire sas_m687;
    reg [63:0] spc687_phy_pc_w;

    

    reg spc688_inst_done;
    wire [1:0]   spc688_thread_id;
    wire [63:0]      spc688_rtl_pc;
    wire sas_m688;
    reg [63:0] spc688_phy_pc_w;

    

    reg spc689_inst_done;
    wire [1:0]   spc689_thread_id;
    wire [63:0]      spc689_rtl_pc;
    wire sas_m689;
    reg [63:0] spc689_phy_pc_w;

    

    reg spc690_inst_done;
    wire [1:0]   spc690_thread_id;
    wire [63:0]      spc690_rtl_pc;
    wire sas_m690;
    reg [63:0] spc690_phy_pc_w;

    

    reg spc691_inst_done;
    wire [1:0]   spc691_thread_id;
    wire [63:0]      spc691_rtl_pc;
    wire sas_m691;
    reg [63:0] spc691_phy_pc_w;

    

    reg spc692_inst_done;
    wire [1:0]   spc692_thread_id;
    wire [63:0]      spc692_rtl_pc;
    wire sas_m692;
    reg [63:0] spc692_phy_pc_w;

    

    reg spc693_inst_done;
    wire [1:0]   spc693_thread_id;
    wire [63:0]      spc693_rtl_pc;
    wire sas_m693;
    reg [63:0] spc693_phy_pc_w;

    

    reg spc694_inst_done;
    wire [1:0]   spc694_thread_id;
    wire [63:0]      spc694_rtl_pc;
    wire sas_m694;
    reg [63:0] spc694_phy_pc_w;

    

    reg spc695_inst_done;
    wire [1:0]   spc695_thread_id;
    wire [63:0]      spc695_rtl_pc;
    wire sas_m695;
    reg [63:0] spc695_phy_pc_w;

    

    reg spc696_inst_done;
    wire [1:0]   spc696_thread_id;
    wire [63:0]      spc696_rtl_pc;
    wire sas_m696;
    reg [63:0] spc696_phy_pc_w;

    

    reg spc697_inst_done;
    wire [1:0]   spc697_thread_id;
    wire [63:0]      spc697_rtl_pc;
    wire sas_m697;
    reg [63:0] spc697_phy_pc_w;

    

    reg spc698_inst_done;
    wire [1:0]   spc698_thread_id;
    wire [63:0]      spc698_rtl_pc;
    wire sas_m698;
    reg [63:0] spc698_phy_pc_w;

    

    reg spc699_inst_done;
    wire [1:0]   spc699_thread_id;
    wire [63:0]      spc699_rtl_pc;
    wire sas_m699;
    reg [63:0] spc699_phy_pc_w;

    

    reg spc700_inst_done;
    wire [1:0]   spc700_thread_id;
    wire [63:0]      spc700_rtl_pc;
    wire sas_m700;
    reg [63:0] spc700_phy_pc_w;

    

    reg spc701_inst_done;
    wire [1:0]   spc701_thread_id;
    wire [63:0]      spc701_rtl_pc;
    wire sas_m701;
    reg [63:0] spc701_phy_pc_w;

    

    reg spc702_inst_done;
    wire [1:0]   spc702_thread_id;
    wire [63:0]      spc702_rtl_pc;
    wire sas_m702;
    reg [63:0] spc702_phy_pc_w;

    

    reg spc703_inst_done;
    wire [1:0]   spc703_thread_id;
    wire [63:0]      spc703_rtl_pc;
    wire sas_m703;
    reg [63:0] spc703_phy_pc_w;

    

    reg spc704_inst_done;
    wire [1:0]   spc704_thread_id;
    wire [63:0]      spc704_rtl_pc;
    wire sas_m704;
    reg [63:0] spc704_phy_pc_w;

    

    reg spc705_inst_done;
    wire [1:0]   spc705_thread_id;
    wire [63:0]      spc705_rtl_pc;
    wire sas_m705;
    reg [63:0] spc705_phy_pc_w;

    

    reg spc706_inst_done;
    wire [1:0]   spc706_thread_id;
    wire [63:0]      spc706_rtl_pc;
    wire sas_m706;
    reg [63:0] spc706_phy_pc_w;

    

    reg spc707_inst_done;
    wire [1:0]   spc707_thread_id;
    wire [63:0]      spc707_rtl_pc;
    wire sas_m707;
    reg [63:0] spc707_phy_pc_w;

    

    reg spc708_inst_done;
    wire [1:0]   spc708_thread_id;
    wire [63:0]      spc708_rtl_pc;
    wire sas_m708;
    reg [63:0] spc708_phy_pc_w;

    

    reg spc709_inst_done;
    wire [1:0]   spc709_thread_id;
    wire [63:0]      spc709_rtl_pc;
    wire sas_m709;
    reg [63:0] spc709_phy_pc_w;

    

    reg spc710_inst_done;
    wire [1:0]   spc710_thread_id;
    wire [63:0]      spc710_rtl_pc;
    wire sas_m710;
    reg [63:0] spc710_phy_pc_w;

    

    reg spc711_inst_done;
    wire [1:0]   spc711_thread_id;
    wire [63:0]      spc711_rtl_pc;
    wire sas_m711;
    reg [63:0] spc711_phy_pc_w;

    

    reg spc712_inst_done;
    wire [1:0]   spc712_thread_id;
    wire [63:0]      spc712_rtl_pc;
    wire sas_m712;
    reg [63:0] spc712_phy_pc_w;

    

    reg spc713_inst_done;
    wire [1:0]   spc713_thread_id;
    wire [63:0]      spc713_rtl_pc;
    wire sas_m713;
    reg [63:0] spc713_phy_pc_w;

    

    reg spc714_inst_done;
    wire [1:0]   spc714_thread_id;
    wire [63:0]      spc714_rtl_pc;
    wire sas_m714;
    reg [63:0] spc714_phy_pc_w;

    

    reg spc715_inst_done;
    wire [1:0]   spc715_thread_id;
    wire [63:0]      spc715_rtl_pc;
    wire sas_m715;
    reg [63:0] spc715_phy_pc_w;

    

    reg spc716_inst_done;
    wire [1:0]   spc716_thread_id;
    wire [63:0]      spc716_rtl_pc;
    wire sas_m716;
    reg [63:0] spc716_phy_pc_w;

    

    reg spc717_inst_done;
    wire [1:0]   spc717_thread_id;
    wire [63:0]      spc717_rtl_pc;
    wire sas_m717;
    reg [63:0] spc717_phy_pc_w;

    

    reg spc718_inst_done;
    wire [1:0]   spc718_thread_id;
    wire [63:0]      spc718_rtl_pc;
    wire sas_m718;
    reg [63:0] spc718_phy_pc_w;

    

    reg spc719_inst_done;
    wire [1:0]   spc719_thread_id;
    wire [63:0]      spc719_rtl_pc;
    wire sas_m719;
    reg [63:0] spc719_phy_pc_w;

    

    reg spc720_inst_done;
    wire [1:0]   spc720_thread_id;
    wire [63:0]      spc720_rtl_pc;
    wire sas_m720;
    reg [63:0] spc720_phy_pc_w;

    

    reg spc721_inst_done;
    wire [1:0]   spc721_thread_id;
    wire [63:0]      spc721_rtl_pc;
    wire sas_m721;
    reg [63:0] spc721_phy_pc_w;

    

    reg spc722_inst_done;
    wire [1:0]   spc722_thread_id;
    wire [63:0]      spc722_rtl_pc;
    wire sas_m722;
    reg [63:0] spc722_phy_pc_w;

    

    reg spc723_inst_done;
    wire [1:0]   spc723_thread_id;
    wire [63:0]      spc723_rtl_pc;
    wire sas_m723;
    reg [63:0] spc723_phy_pc_w;

    

    reg spc724_inst_done;
    wire [1:0]   spc724_thread_id;
    wire [63:0]      spc724_rtl_pc;
    wire sas_m724;
    reg [63:0] spc724_phy_pc_w;

    

    reg spc725_inst_done;
    wire [1:0]   spc725_thread_id;
    wire [63:0]      spc725_rtl_pc;
    wire sas_m725;
    reg [63:0] spc725_phy_pc_w;

    

    reg spc726_inst_done;
    wire [1:0]   spc726_thread_id;
    wire [63:0]      spc726_rtl_pc;
    wire sas_m726;
    reg [63:0] spc726_phy_pc_w;

    

    reg spc727_inst_done;
    wire [1:0]   spc727_thread_id;
    wire [63:0]      spc727_rtl_pc;
    wire sas_m727;
    reg [63:0] spc727_phy_pc_w;

    

    reg spc728_inst_done;
    wire [1:0]   spc728_thread_id;
    wire [63:0]      spc728_rtl_pc;
    wire sas_m728;
    reg [63:0] spc728_phy_pc_w;

    

    reg spc729_inst_done;
    wire [1:0]   spc729_thread_id;
    wire [63:0]      spc729_rtl_pc;
    wire sas_m729;
    reg [63:0] spc729_phy_pc_w;

    

    reg spc730_inst_done;
    wire [1:0]   spc730_thread_id;
    wire [63:0]      spc730_rtl_pc;
    wire sas_m730;
    reg [63:0] spc730_phy_pc_w;

    

    reg spc731_inst_done;
    wire [1:0]   spc731_thread_id;
    wire [63:0]      spc731_rtl_pc;
    wire sas_m731;
    reg [63:0] spc731_phy_pc_w;

    

    reg spc732_inst_done;
    wire [1:0]   spc732_thread_id;
    wire [63:0]      spc732_rtl_pc;
    wire sas_m732;
    reg [63:0] spc732_phy_pc_w;

    

    reg spc733_inst_done;
    wire [1:0]   spc733_thread_id;
    wire [63:0]      spc733_rtl_pc;
    wire sas_m733;
    reg [63:0] spc733_phy_pc_w;

    

    reg spc734_inst_done;
    wire [1:0]   spc734_thread_id;
    wire [63:0]      spc734_rtl_pc;
    wire sas_m734;
    reg [63:0] spc734_phy_pc_w;

    

    reg spc735_inst_done;
    wire [1:0]   spc735_thread_id;
    wire [63:0]      spc735_rtl_pc;
    wire sas_m735;
    reg [63:0] spc735_phy_pc_w;

    

    reg spc736_inst_done;
    wire [1:0]   spc736_thread_id;
    wire [63:0]      spc736_rtl_pc;
    wire sas_m736;
    reg [63:0] spc736_phy_pc_w;

    

    reg spc737_inst_done;
    wire [1:0]   spc737_thread_id;
    wire [63:0]      spc737_rtl_pc;
    wire sas_m737;
    reg [63:0] spc737_phy_pc_w;

    

    reg spc738_inst_done;
    wire [1:0]   spc738_thread_id;
    wire [63:0]      spc738_rtl_pc;
    wire sas_m738;
    reg [63:0] spc738_phy_pc_w;

    

    reg spc739_inst_done;
    wire [1:0]   spc739_thread_id;
    wire [63:0]      spc739_rtl_pc;
    wire sas_m739;
    reg [63:0] spc739_phy_pc_w;

    

    reg spc740_inst_done;
    wire [1:0]   spc740_thread_id;
    wire [63:0]      spc740_rtl_pc;
    wire sas_m740;
    reg [63:0] spc740_phy_pc_w;

    

    reg spc741_inst_done;
    wire [1:0]   spc741_thread_id;
    wire [63:0]      spc741_rtl_pc;
    wire sas_m741;
    reg [63:0] spc741_phy_pc_w;

    

    reg spc742_inst_done;
    wire [1:0]   spc742_thread_id;
    wire [63:0]      spc742_rtl_pc;
    wire sas_m742;
    reg [63:0] spc742_phy_pc_w;

    

    reg spc743_inst_done;
    wire [1:0]   spc743_thread_id;
    wire [63:0]      spc743_rtl_pc;
    wire sas_m743;
    reg [63:0] spc743_phy_pc_w;

    

    reg spc744_inst_done;
    wire [1:0]   spc744_thread_id;
    wire [63:0]      spc744_rtl_pc;
    wire sas_m744;
    reg [63:0] spc744_phy_pc_w;

    

    reg spc745_inst_done;
    wire [1:0]   spc745_thread_id;
    wire [63:0]      spc745_rtl_pc;
    wire sas_m745;
    reg [63:0] spc745_phy_pc_w;

    

    reg spc746_inst_done;
    wire [1:0]   spc746_thread_id;
    wire [63:0]      spc746_rtl_pc;
    wire sas_m746;
    reg [63:0] spc746_phy_pc_w;

    

    reg spc747_inst_done;
    wire [1:0]   spc747_thread_id;
    wire [63:0]      spc747_rtl_pc;
    wire sas_m747;
    reg [63:0] spc747_phy_pc_w;

    

    reg spc748_inst_done;
    wire [1:0]   spc748_thread_id;
    wire [63:0]      spc748_rtl_pc;
    wire sas_m748;
    reg [63:0] spc748_phy_pc_w;

    

    reg spc749_inst_done;
    wire [1:0]   spc749_thread_id;
    wire [63:0]      spc749_rtl_pc;
    wire sas_m749;
    reg [63:0] spc749_phy_pc_w;

    

    reg spc750_inst_done;
    wire [1:0]   spc750_thread_id;
    wire [63:0]      spc750_rtl_pc;
    wire sas_m750;
    reg [63:0] spc750_phy_pc_w;

    

    reg spc751_inst_done;
    wire [1:0]   spc751_thread_id;
    wire [63:0]      spc751_rtl_pc;
    wire sas_m751;
    reg [63:0] spc751_phy_pc_w;

    

    reg spc752_inst_done;
    wire [1:0]   spc752_thread_id;
    wire [63:0]      spc752_rtl_pc;
    wire sas_m752;
    reg [63:0] spc752_phy_pc_w;

    

    reg spc753_inst_done;
    wire [1:0]   spc753_thread_id;
    wire [63:0]      spc753_rtl_pc;
    wire sas_m753;
    reg [63:0] spc753_phy_pc_w;

    

    reg spc754_inst_done;
    wire [1:0]   spc754_thread_id;
    wire [63:0]      spc754_rtl_pc;
    wire sas_m754;
    reg [63:0] spc754_phy_pc_w;

    

    reg spc755_inst_done;
    wire [1:0]   spc755_thread_id;
    wire [63:0]      spc755_rtl_pc;
    wire sas_m755;
    reg [63:0] spc755_phy_pc_w;

    

    reg spc756_inst_done;
    wire [1:0]   spc756_thread_id;
    wire [63:0]      spc756_rtl_pc;
    wire sas_m756;
    reg [63:0] spc756_phy_pc_w;

    

    reg spc757_inst_done;
    wire [1:0]   spc757_thread_id;
    wire [63:0]      spc757_rtl_pc;
    wire sas_m757;
    reg [63:0] spc757_phy_pc_w;

    

    reg spc758_inst_done;
    wire [1:0]   spc758_thread_id;
    wire [63:0]      spc758_rtl_pc;
    wire sas_m758;
    reg [63:0] spc758_phy_pc_w;

    

    reg spc759_inst_done;
    wire [1:0]   spc759_thread_id;
    wire [63:0]      spc759_rtl_pc;
    wire sas_m759;
    reg [63:0] spc759_phy_pc_w;

    

    reg spc760_inst_done;
    wire [1:0]   spc760_thread_id;
    wire [63:0]      spc760_rtl_pc;
    wire sas_m760;
    reg [63:0] spc760_phy_pc_w;

    

    reg spc761_inst_done;
    wire [1:0]   spc761_thread_id;
    wire [63:0]      spc761_rtl_pc;
    wire sas_m761;
    reg [63:0] spc761_phy_pc_w;

    

    reg spc762_inst_done;
    wire [1:0]   spc762_thread_id;
    wire [63:0]      spc762_rtl_pc;
    wire sas_m762;
    reg [63:0] spc762_phy_pc_w;

    

    reg spc763_inst_done;
    wire [1:0]   spc763_thread_id;
    wire [63:0]      spc763_rtl_pc;
    wire sas_m763;
    reg [63:0] spc763_phy_pc_w;

    

    reg spc764_inst_done;
    wire [1:0]   spc764_thread_id;
    wire [63:0]      spc764_rtl_pc;
    wire sas_m764;
    reg [63:0] spc764_phy_pc_w;

    

    reg spc765_inst_done;
    wire [1:0]   spc765_thread_id;
    wire [63:0]      spc765_rtl_pc;
    wire sas_m765;
    reg [63:0] spc765_phy_pc_w;

    

    reg spc766_inst_done;
    wire [1:0]   spc766_thread_id;
    wire [63:0]      spc766_rtl_pc;
    wire sas_m766;
    reg [63:0] spc766_phy_pc_w;

    

    reg spc767_inst_done;
    wire [1:0]   spc767_thread_id;
    wire [63:0]      spc767_rtl_pc;
    wire sas_m767;
    reg [63:0] spc767_phy_pc_w;

    

    reg spc768_inst_done;
    wire [1:0]   spc768_thread_id;
    wire [63:0]      spc768_rtl_pc;
    wire sas_m768;
    reg [63:0] spc768_phy_pc_w;

    

    reg spc769_inst_done;
    wire [1:0]   spc769_thread_id;
    wire [63:0]      spc769_rtl_pc;
    wire sas_m769;
    reg [63:0] spc769_phy_pc_w;

    

    reg spc770_inst_done;
    wire [1:0]   spc770_thread_id;
    wire [63:0]      spc770_rtl_pc;
    wire sas_m770;
    reg [63:0] spc770_phy_pc_w;

    

    reg spc771_inst_done;
    wire [1:0]   spc771_thread_id;
    wire [63:0]      spc771_rtl_pc;
    wire sas_m771;
    reg [63:0] spc771_phy_pc_w;

    

    reg spc772_inst_done;
    wire [1:0]   spc772_thread_id;
    wire [63:0]      spc772_rtl_pc;
    wire sas_m772;
    reg [63:0] spc772_phy_pc_w;

    

    reg spc773_inst_done;
    wire [1:0]   spc773_thread_id;
    wire [63:0]      spc773_rtl_pc;
    wire sas_m773;
    reg [63:0] spc773_phy_pc_w;

    

    reg spc774_inst_done;
    wire [1:0]   spc774_thread_id;
    wire [63:0]      spc774_rtl_pc;
    wire sas_m774;
    reg [63:0] spc774_phy_pc_w;

    

    reg spc775_inst_done;
    wire [1:0]   spc775_thread_id;
    wire [63:0]      spc775_rtl_pc;
    wire sas_m775;
    reg [63:0] spc775_phy_pc_w;

    

    reg spc776_inst_done;
    wire [1:0]   spc776_thread_id;
    wire [63:0]      spc776_rtl_pc;
    wire sas_m776;
    reg [63:0] spc776_phy_pc_w;

    

    reg spc777_inst_done;
    wire [1:0]   spc777_thread_id;
    wire [63:0]      spc777_rtl_pc;
    wire sas_m777;
    reg [63:0] spc777_phy_pc_w;

    

    reg spc778_inst_done;
    wire [1:0]   spc778_thread_id;
    wire [63:0]      spc778_rtl_pc;
    wire sas_m778;
    reg [63:0] spc778_phy_pc_w;

    

    reg spc779_inst_done;
    wire [1:0]   spc779_thread_id;
    wire [63:0]      spc779_rtl_pc;
    wire sas_m779;
    reg [63:0] spc779_phy_pc_w;

    

    reg spc780_inst_done;
    wire [1:0]   spc780_thread_id;
    wire [63:0]      spc780_rtl_pc;
    wire sas_m780;
    reg [63:0] spc780_phy_pc_w;

    

    reg spc781_inst_done;
    wire [1:0]   spc781_thread_id;
    wire [63:0]      spc781_rtl_pc;
    wire sas_m781;
    reg [63:0] spc781_phy_pc_w;

    

    reg spc782_inst_done;
    wire [1:0]   spc782_thread_id;
    wire [63:0]      spc782_rtl_pc;
    wire sas_m782;
    reg [63:0] spc782_phy_pc_w;

    

    reg spc783_inst_done;
    wire [1:0]   spc783_thread_id;
    wire [63:0]      spc783_rtl_pc;
    wire sas_m783;
    reg [63:0] spc783_phy_pc_w;

    

    reg spc784_inst_done;
    wire [1:0]   spc784_thread_id;
    wire [63:0]      spc784_rtl_pc;
    wire sas_m784;
    reg [63:0] spc784_phy_pc_w;

    

    reg spc785_inst_done;
    wire [1:0]   spc785_thread_id;
    wire [63:0]      spc785_rtl_pc;
    wire sas_m785;
    reg [63:0] spc785_phy_pc_w;

    

    reg spc786_inst_done;
    wire [1:0]   spc786_thread_id;
    wire [63:0]      spc786_rtl_pc;
    wire sas_m786;
    reg [63:0] spc786_phy_pc_w;

    

    reg spc787_inst_done;
    wire [1:0]   spc787_thread_id;
    wire [63:0]      spc787_rtl_pc;
    wire sas_m787;
    reg [63:0] spc787_phy_pc_w;

    

    reg spc788_inst_done;
    wire [1:0]   spc788_thread_id;
    wire [63:0]      spc788_rtl_pc;
    wire sas_m788;
    reg [63:0] spc788_phy_pc_w;

    

    reg spc789_inst_done;
    wire [1:0]   spc789_thread_id;
    wire [63:0]      spc789_rtl_pc;
    wire sas_m789;
    reg [63:0] spc789_phy_pc_w;

    

    reg spc790_inst_done;
    wire [1:0]   spc790_thread_id;
    wire [63:0]      spc790_rtl_pc;
    wire sas_m790;
    reg [63:0] spc790_phy_pc_w;

    

    reg spc791_inst_done;
    wire [1:0]   spc791_thread_id;
    wire [63:0]      spc791_rtl_pc;
    wire sas_m791;
    reg [63:0] spc791_phy_pc_w;

    

    reg spc792_inst_done;
    wire [1:0]   spc792_thread_id;
    wire [63:0]      spc792_rtl_pc;
    wire sas_m792;
    reg [63:0] spc792_phy_pc_w;

    

    reg spc793_inst_done;
    wire [1:0]   spc793_thread_id;
    wire [63:0]      spc793_rtl_pc;
    wire sas_m793;
    reg [63:0] spc793_phy_pc_w;

    

    reg spc794_inst_done;
    wire [1:0]   spc794_thread_id;
    wire [63:0]      spc794_rtl_pc;
    wire sas_m794;
    reg [63:0] spc794_phy_pc_w;

    

    reg spc795_inst_done;
    wire [1:0]   spc795_thread_id;
    wire [63:0]      spc795_rtl_pc;
    wire sas_m795;
    reg [63:0] spc795_phy_pc_w;

    

    reg spc796_inst_done;
    wire [1:0]   spc796_thread_id;
    wire [63:0]      spc796_rtl_pc;
    wire sas_m796;
    reg [63:0] spc796_phy_pc_w;

    

    reg spc797_inst_done;
    wire [1:0]   spc797_thread_id;
    wire [63:0]      spc797_rtl_pc;
    wire sas_m797;
    reg [63:0] spc797_phy_pc_w;

    

    reg spc798_inst_done;
    wire [1:0]   spc798_thread_id;
    wire [63:0]      spc798_rtl_pc;
    wire sas_m798;
    reg [63:0] spc798_phy_pc_w;

    

    reg spc799_inst_done;
    wire [1:0]   spc799_thread_id;
    wire [63:0]      spc799_rtl_pc;
    wire sas_m799;
    reg [63:0] spc799_phy_pc_w;

    

    reg spc800_inst_done;
    wire [1:0]   spc800_thread_id;
    wire [63:0]      spc800_rtl_pc;
    wire sas_m800;
    reg [63:0] spc800_phy_pc_w;

    

    reg spc801_inst_done;
    wire [1:0]   spc801_thread_id;
    wire [63:0]      spc801_rtl_pc;
    wire sas_m801;
    reg [63:0] spc801_phy_pc_w;

    

    reg spc802_inst_done;
    wire [1:0]   spc802_thread_id;
    wire [63:0]      spc802_rtl_pc;
    wire sas_m802;
    reg [63:0] spc802_phy_pc_w;

    

    reg spc803_inst_done;
    wire [1:0]   spc803_thread_id;
    wire [63:0]      spc803_rtl_pc;
    wire sas_m803;
    reg [63:0] spc803_phy_pc_w;

    

    reg spc804_inst_done;
    wire [1:0]   spc804_thread_id;
    wire [63:0]      spc804_rtl_pc;
    wire sas_m804;
    reg [63:0] spc804_phy_pc_w;

    

    reg spc805_inst_done;
    wire [1:0]   spc805_thread_id;
    wire [63:0]      spc805_rtl_pc;
    wire sas_m805;
    reg [63:0] spc805_phy_pc_w;

    

    reg spc806_inst_done;
    wire [1:0]   spc806_thread_id;
    wire [63:0]      spc806_rtl_pc;
    wire sas_m806;
    reg [63:0] spc806_phy_pc_w;

    

    reg spc807_inst_done;
    wire [1:0]   spc807_thread_id;
    wire [63:0]      spc807_rtl_pc;
    wire sas_m807;
    reg [63:0] spc807_phy_pc_w;

    

    reg spc808_inst_done;
    wire [1:0]   spc808_thread_id;
    wire [63:0]      spc808_rtl_pc;
    wire sas_m808;
    reg [63:0] spc808_phy_pc_w;

    

    reg spc809_inst_done;
    wire [1:0]   spc809_thread_id;
    wire [63:0]      spc809_rtl_pc;
    wire sas_m809;
    reg [63:0] spc809_phy_pc_w;

    

    reg spc810_inst_done;
    wire [1:0]   spc810_thread_id;
    wire [63:0]      spc810_rtl_pc;
    wire sas_m810;
    reg [63:0] spc810_phy_pc_w;

    

    reg spc811_inst_done;
    wire [1:0]   spc811_thread_id;
    wire [63:0]      spc811_rtl_pc;
    wire sas_m811;
    reg [63:0] spc811_phy_pc_w;

    

    reg spc812_inst_done;
    wire [1:0]   spc812_thread_id;
    wire [63:0]      spc812_rtl_pc;
    wire sas_m812;
    reg [63:0] spc812_phy_pc_w;

    

    reg spc813_inst_done;
    wire [1:0]   spc813_thread_id;
    wire [63:0]      spc813_rtl_pc;
    wire sas_m813;
    reg [63:0] spc813_phy_pc_w;

    

    reg spc814_inst_done;
    wire [1:0]   spc814_thread_id;
    wire [63:0]      spc814_rtl_pc;
    wire sas_m814;
    reg [63:0] spc814_phy_pc_w;

    

    reg spc815_inst_done;
    wire [1:0]   spc815_thread_id;
    wire [63:0]      spc815_rtl_pc;
    wire sas_m815;
    reg [63:0] spc815_phy_pc_w;

    

    reg spc816_inst_done;
    wire [1:0]   spc816_thread_id;
    wire [63:0]      spc816_rtl_pc;
    wire sas_m816;
    reg [63:0] spc816_phy_pc_w;

    

    reg spc817_inst_done;
    wire [1:0]   spc817_thread_id;
    wire [63:0]      spc817_rtl_pc;
    wire sas_m817;
    reg [63:0] spc817_phy_pc_w;

    

    reg spc818_inst_done;
    wire [1:0]   spc818_thread_id;
    wire [63:0]      spc818_rtl_pc;
    wire sas_m818;
    reg [63:0] spc818_phy_pc_w;

    

    reg spc819_inst_done;
    wire [1:0]   spc819_thread_id;
    wire [63:0]      spc819_rtl_pc;
    wire sas_m819;
    reg [63:0] spc819_phy_pc_w;

    

    reg spc820_inst_done;
    wire [1:0]   spc820_thread_id;
    wire [63:0]      spc820_rtl_pc;
    wire sas_m820;
    reg [63:0] spc820_phy_pc_w;

    

    reg spc821_inst_done;
    wire [1:0]   spc821_thread_id;
    wire [63:0]      spc821_rtl_pc;
    wire sas_m821;
    reg [63:0] spc821_phy_pc_w;

    

    reg spc822_inst_done;
    wire [1:0]   spc822_thread_id;
    wire [63:0]      spc822_rtl_pc;
    wire sas_m822;
    reg [63:0] spc822_phy_pc_w;

    

    reg spc823_inst_done;
    wire [1:0]   spc823_thread_id;
    wire [63:0]      spc823_rtl_pc;
    wire sas_m823;
    reg [63:0] spc823_phy_pc_w;

    

    reg spc824_inst_done;
    wire [1:0]   spc824_thread_id;
    wire [63:0]      spc824_rtl_pc;
    wire sas_m824;
    reg [63:0] spc824_phy_pc_w;

    

    reg spc825_inst_done;
    wire [1:0]   spc825_thread_id;
    wire [63:0]      spc825_rtl_pc;
    wire sas_m825;
    reg [63:0] spc825_phy_pc_w;

    

    reg spc826_inst_done;
    wire [1:0]   spc826_thread_id;
    wire [63:0]      spc826_rtl_pc;
    wire sas_m826;
    reg [63:0] spc826_phy_pc_w;

    

    reg spc827_inst_done;
    wire [1:0]   spc827_thread_id;
    wire [63:0]      spc827_rtl_pc;
    wire sas_m827;
    reg [63:0] spc827_phy_pc_w;

    

    reg spc828_inst_done;
    wire [1:0]   spc828_thread_id;
    wire [63:0]      spc828_rtl_pc;
    wire sas_m828;
    reg [63:0] spc828_phy_pc_w;

    

    reg spc829_inst_done;
    wire [1:0]   spc829_thread_id;
    wire [63:0]      spc829_rtl_pc;
    wire sas_m829;
    reg [63:0] spc829_phy_pc_w;

    

    reg spc830_inst_done;
    wire [1:0]   spc830_thread_id;
    wire [63:0]      spc830_rtl_pc;
    wire sas_m830;
    reg [63:0] spc830_phy_pc_w;

    

    reg spc831_inst_done;
    wire [1:0]   spc831_thread_id;
    wire [63:0]      spc831_rtl_pc;
    wire sas_m831;
    reg [63:0] spc831_phy_pc_w;

    

    reg spc832_inst_done;
    wire [1:0]   spc832_thread_id;
    wire [63:0]      spc832_rtl_pc;
    wire sas_m832;
    reg [63:0] spc832_phy_pc_w;

    

    reg spc833_inst_done;
    wire [1:0]   spc833_thread_id;
    wire [63:0]      spc833_rtl_pc;
    wire sas_m833;
    reg [63:0] spc833_phy_pc_w;

    

    reg spc834_inst_done;
    wire [1:0]   spc834_thread_id;
    wire [63:0]      spc834_rtl_pc;
    wire sas_m834;
    reg [63:0] spc834_phy_pc_w;

    

    reg spc835_inst_done;
    wire [1:0]   spc835_thread_id;
    wire [63:0]      spc835_rtl_pc;
    wire sas_m835;
    reg [63:0] spc835_phy_pc_w;

    

    reg spc836_inst_done;
    wire [1:0]   spc836_thread_id;
    wire [63:0]      spc836_rtl_pc;
    wire sas_m836;
    reg [63:0] spc836_phy_pc_w;

    

    reg spc837_inst_done;
    wire [1:0]   spc837_thread_id;
    wire [63:0]      spc837_rtl_pc;
    wire sas_m837;
    reg [63:0] spc837_phy_pc_w;

    

    reg spc838_inst_done;
    wire [1:0]   spc838_thread_id;
    wire [63:0]      spc838_rtl_pc;
    wire sas_m838;
    reg [63:0] spc838_phy_pc_w;

    

    reg spc839_inst_done;
    wire [1:0]   spc839_thread_id;
    wire [63:0]      spc839_rtl_pc;
    wire sas_m839;
    reg [63:0] spc839_phy_pc_w;

    

    reg spc840_inst_done;
    wire [1:0]   spc840_thread_id;
    wire [63:0]      spc840_rtl_pc;
    wire sas_m840;
    reg [63:0] spc840_phy_pc_w;

    

    reg spc841_inst_done;
    wire [1:0]   spc841_thread_id;
    wire [63:0]      spc841_rtl_pc;
    wire sas_m841;
    reg [63:0] spc841_phy_pc_w;

    

    reg spc842_inst_done;
    wire [1:0]   spc842_thread_id;
    wire [63:0]      spc842_rtl_pc;
    wire sas_m842;
    reg [63:0] spc842_phy_pc_w;

    

    reg spc843_inst_done;
    wire [1:0]   spc843_thread_id;
    wire [63:0]      spc843_rtl_pc;
    wire sas_m843;
    reg [63:0] spc843_phy_pc_w;

    

    reg spc844_inst_done;
    wire [1:0]   spc844_thread_id;
    wire [63:0]      spc844_rtl_pc;
    wire sas_m844;
    reg [63:0] spc844_phy_pc_w;

    

    reg spc845_inst_done;
    wire [1:0]   spc845_thread_id;
    wire [63:0]      spc845_rtl_pc;
    wire sas_m845;
    reg [63:0] spc845_phy_pc_w;

    

    reg spc846_inst_done;
    wire [1:0]   spc846_thread_id;
    wire [63:0]      spc846_rtl_pc;
    wire sas_m846;
    reg [63:0] spc846_phy_pc_w;

    

    reg spc847_inst_done;
    wire [1:0]   spc847_thread_id;
    wire [63:0]      spc847_rtl_pc;
    wire sas_m847;
    reg [63:0] spc847_phy_pc_w;

    

    reg spc848_inst_done;
    wire [1:0]   spc848_thread_id;
    wire [63:0]      spc848_rtl_pc;
    wire sas_m848;
    reg [63:0] spc848_phy_pc_w;

    

    reg spc849_inst_done;
    wire [1:0]   spc849_thread_id;
    wire [63:0]      spc849_rtl_pc;
    wire sas_m849;
    reg [63:0] spc849_phy_pc_w;

    

    reg spc850_inst_done;
    wire [1:0]   spc850_thread_id;
    wire [63:0]      spc850_rtl_pc;
    wire sas_m850;
    reg [63:0] spc850_phy_pc_w;

    

    reg spc851_inst_done;
    wire [1:0]   spc851_thread_id;
    wire [63:0]      spc851_rtl_pc;
    wire sas_m851;
    reg [63:0] spc851_phy_pc_w;

    

    reg spc852_inst_done;
    wire [1:0]   spc852_thread_id;
    wire [63:0]      spc852_rtl_pc;
    wire sas_m852;
    reg [63:0] spc852_phy_pc_w;

    

    reg spc853_inst_done;
    wire [1:0]   spc853_thread_id;
    wire [63:0]      spc853_rtl_pc;
    wire sas_m853;
    reg [63:0] spc853_phy_pc_w;

    

    reg spc854_inst_done;
    wire [1:0]   spc854_thread_id;
    wire [63:0]      spc854_rtl_pc;
    wire sas_m854;
    reg [63:0] spc854_phy_pc_w;

    

    reg spc855_inst_done;
    wire [1:0]   spc855_thread_id;
    wire [63:0]      spc855_rtl_pc;
    wire sas_m855;
    reg [63:0] spc855_phy_pc_w;

    

    reg spc856_inst_done;
    wire [1:0]   spc856_thread_id;
    wire [63:0]      spc856_rtl_pc;
    wire sas_m856;
    reg [63:0] spc856_phy_pc_w;

    

    reg spc857_inst_done;
    wire [1:0]   spc857_thread_id;
    wire [63:0]      spc857_rtl_pc;
    wire sas_m857;
    reg [63:0] spc857_phy_pc_w;

    

    reg spc858_inst_done;
    wire [1:0]   spc858_thread_id;
    wire [63:0]      spc858_rtl_pc;
    wire sas_m858;
    reg [63:0] spc858_phy_pc_w;

    

    reg spc859_inst_done;
    wire [1:0]   spc859_thread_id;
    wire [63:0]      spc859_rtl_pc;
    wire sas_m859;
    reg [63:0] spc859_phy_pc_w;

    

    reg spc860_inst_done;
    wire [1:0]   spc860_thread_id;
    wire [63:0]      spc860_rtl_pc;
    wire sas_m860;
    reg [63:0] spc860_phy_pc_w;

    

    reg spc861_inst_done;
    wire [1:0]   spc861_thread_id;
    wire [63:0]      spc861_rtl_pc;
    wire sas_m861;
    reg [63:0] spc861_phy_pc_w;

    

    reg spc862_inst_done;
    wire [1:0]   spc862_thread_id;
    wire [63:0]      spc862_rtl_pc;
    wire sas_m862;
    reg [63:0] spc862_phy_pc_w;

    

    reg spc863_inst_done;
    wire [1:0]   spc863_thread_id;
    wire [63:0]      spc863_rtl_pc;
    wire sas_m863;
    reg [63:0] spc863_phy_pc_w;

    

    reg spc864_inst_done;
    wire [1:0]   spc864_thread_id;
    wire [63:0]      spc864_rtl_pc;
    wire sas_m864;
    reg [63:0] spc864_phy_pc_w;

    

    reg spc865_inst_done;
    wire [1:0]   spc865_thread_id;
    wire [63:0]      spc865_rtl_pc;
    wire sas_m865;
    reg [63:0] spc865_phy_pc_w;

    

    reg spc866_inst_done;
    wire [1:0]   spc866_thread_id;
    wire [63:0]      spc866_rtl_pc;
    wire sas_m866;
    reg [63:0] spc866_phy_pc_w;

    

    reg spc867_inst_done;
    wire [1:0]   spc867_thread_id;
    wire [63:0]      spc867_rtl_pc;
    wire sas_m867;
    reg [63:0] spc867_phy_pc_w;

    

    reg spc868_inst_done;
    wire [1:0]   spc868_thread_id;
    wire [63:0]      spc868_rtl_pc;
    wire sas_m868;
    reg [63:0] spc868_phy_pc_w;

    

    reg spc869_inst_done;
    wire [1:0]   spc869_thread_id;
    wire [63:0]      spc869_rtl_pc;
    wire sas_m869;
    reg [63:0] spc869_phy_pc_w;

    

    reg spc870_inst_done;
    wire [1:0]   spc870_thread_id;
    wire [63:0]      spc870_rtl_pc;
    wire sas_m870;
    reg [63:0] spc870_phy_pc_w;

    

    reg spc871_inst_done;
    wire [1:0]   spc871_thread_id;
    wire [63:0]      spc871_rtl_pc;
    wire sas_m871;
    reg [63:0] spc871_phy_pc_w;

    

    reg spc872_inst_done;
    wire [1:0]   spc872_thread_id;
    wire [63:0]      spc872_rtl_pc;
    wire sas_m872;
    reg [63:0] spc872_phy_pc_w;

    

    reg spc873_inst_done;
    wire [1:0]   spc873_thread_id;
    wire [63:0]      spc873_rtl_pc;
    wire sas_m873;
    reg [63:0] spc873_phy_pc_w;

    

    reg spc874_inst_done;
    wire [1:0]   spc874_thread_id;
    wire [63:0]      spc874_rtl_pc;
    wire sas_m874;
    reg [63:0] spc874_phy_pc_w;

    

    reg spc875_inst_done;
    wire [1:0]   spc875_thread_id;
    wire [63:0]      spc875_rtl_pc;
    wire sas_m875;
    reg [63:0] spc875_phy_pc_w;

    

    reg spc876_inst_done;
    wire [1:0]   spc876_thread_id;
    wire [63:0]      spc876_rtl_pc;
    wire sas_m876;
    reg [63:0] spc876_phy_pc_w;

    

    reg spc877_inst_done;
    wire [1:0]   spc877_thread_id;
    wire [63:0]      spc877_rtl_pc;
    wire sas_m877;
    reg [63:0] spc877_phy_pc_w;

    

    reg spc878_inst_done;
    wire [1:0]   spc878_thread_id;
    wire [63:0]      spc878_rtl_pc;
    wire sas_m878;
    reg [63:0] spc878_phy_pc_w;

    

    reg spc879_inst_done;
    wire [1:0]   spc879_thread_id;
    wire [63:0]      spc879_rtl_pc;
    wire sas_m879;
    reg [63:0] spc879_phy_pc_w;

    

    reg spc880_inst_done;
    wire [1:0]   spc880_thread_id;
    wire [63:0]      spc880_rtl_pc;
    wire sas_m880;
    reg [63:0] spc880_phy_pc_w;

    

    reg spc881_inst_done;
    wire [1:0]   spc881_thread_id;
    wire [63:0]      spc881_rtl_pc;
    wire sas_m881;
    reg [63:0] spc881_phy_pc_w;

    

    reg spc882_inst_done;
    wire [1:0]   spc882_thread_id;
    wire [63:0]      spc882_rtl_pc;
    wire sas_m882;
    reg [63:0] spc882_phy_pc_w;

    

    reg spc883_inst_done;
    wire [1:0]   spc883_thread_id;
    wire [63:0]      spc883_rtl_pc;
    wire sas_m883;
    reg [63:0] spc883_phy_pc_w;

    

    reg spc884_inst_done;
    wire [1:0]   spc884_thread_id;
    wire [63:0]      spc884_rtl_pc;
    wire sas_m884;
    reg [63:0] spc884_phy_pc_w;

    

    reg spc885_inst_done;
    wire [1:0]   spc885_thread_id;
    wire [63:0]      spc885_rtl_pc;
    wire sas_m885;
    reg [63:0] spc885_phy_pc_w;

    

    reg spc886_inst_done;
    wire [1:0]   spc886_thread_id;
    wire [63:0]      spc886_rtl_pc;
    wire sas_m886;
    reg [63:0] spc886_phy_pc_w;

    

    reg spc887_inst_done;
    wire [1:0]   spc887_thread_id;
    wire [63:0]      spc887_rtl_pc;
    wire sas_m887;
    reg [63:0] spc887_phy_pc_w;

    

    reg spc888_inst_done;
    wire [1:0]   spc888_thread_id;
    wire [63:0]      spc888_rtl_pc;
    wire sas_m888;
    reg [63:0] spc888_phy_pc_w;

    

    reg spc889_inst_done;
    wire [1:0]   spc889_thread_id;
    wire [63:0]      spc889_rtl_pc;
    wire sas_m889;
    reg [63:0] spc889_phy_pc_w;

    

    reg spc890_inst_done;
    wire [1:0]   spc890_thread_id;
    wire [63:0]      spc890_rtl_pc;
    wire sas_m890;
    reg [63:0] spc890_phy_pc_w;

    

    reg spc891_inst_done;
    wire [1:0]   spc891_thread_id;
    wire [63:0]      spc891_rtl_pc;
    wire sas_m891;
    reg [63:0] spc891_phy_pc_w;

    

    reg spc892_inst_done;
    wire [1:0]   spc892_thread_id;
    wire [63:0]      spc892_rtl_pc;
    wire sas_m892;
    reg [63:0] spc892_phy_pc_w;

    

    reg spc893_inst_done;
    wire [1:0]   spc893_thread_id;
    wire [63:0]      spc893_rtl_pc;
    wire sas_m893;
    reg [63:0] spc893_phy_pc_w;

    

    reg spc894_inst_done;
    wire [1:0]   spc894_thread_id;
    wire [63:0]      spc894_rtl_pc;
    wire sas_m894;
    reg [63:0] spc894_phy_pc_w;

    

    reg spc895_inst_done;
    wire [1:0]   spc895_thread_id;
    wire [63:0]      spc895_rtl_pc;
    wire sas_m895;
    reg [63:0] spc895_phy_pc_w;

    

    reg spc896_inst_done;
    wire [1:0]   spc896_thread_id;
    wire [63:0]      spc896_rtl_pc;
    wire sas_m896;
    reg [63:0] spc896_phy_pc_w;

    

    reg spc897_inst_done;
    wire [1:0]   spc897_thread_id;
    wire [63:0]      spc897_rtl_pc;
    wire sas_m897;
    reg [63:0] spc897_phy_pc_w;

    

    reg spc898_inst_done;
    wire [1:0]   spc898_thread_id;
    wire [63:0]      spc898_rtl_pc;
    wire sas_m898;
    reg [63:0] spc898_phy_pc_w;

    

    reg spc899_inst_done;
    wire [1:0]   spc899_thread_id;
    wire [63:0]      spc899_rtl_pc;
    wire sas_m899;
    reg [63:0] spc899_phy_pc_w;

    

    reg spc900_inst_done;
    wire [1:0]   spc900_thread_id;
    wire [63:0]      spc900_rtl_pc;
    wire sas_m900;
    reg [63:0] spc900_phy_pc_w;

    

    reg spc901_inst_done;
    wire [1:0]   spc901_thread_id;
    wire [63:0]      spc901_rtl_pc;
    wire sas_m901;
    reg [63:0] spc901_phy_pc_w;

    

    reg spc902_inst_done;
    wire [1:0]   spc902_thread_id;
    wire [63:0]      spc902_rtl_pc;
    wire sas_m902;
    reg [63:0] spc902_phy_pc_w;

    

    reg spc903_inst_done;
    wire [1:0]   spc903_thread_id;
    wire [63:0]      spc903_rtl_pc;
    wire sas_m903;
    reg [63:0] spc903_phy_pc_w;

    

    reg spc904_inst_done;
    wire [1:0]   spc904_thread_id;
    wire [63:0]      spc904_rtl_pc;
    wire sas_m904;
    reg [63:0] spc904_phy_pc_w;

    

    reg spc905_inst_done;
    wire [1:0]   spc905_thread_id;
    wire [63:0]      spc905_rtl_pc;
    wire sas_m905;
    reg [63:0] spc905_phy_pc_w;

    

    reg spc906_inst_done;
    wire [1:0]   spc906_thread_id;
    wire [63:0]      spc906_rtl_pc;
    wire sas_m906;
    reg [63:0] spc906_phy_pc_w;

    

    reg spc907_inst_done;
    wire [1:0]   spc907_thread_id;
    wire [63:0]      spc907_rtl_pc;
    wire sas_m907;
    reg [63:0] spc907_phy_pc_w;

    

    reg spc908_inst_done;
    wire [1:0]   spc908_thread_id;
    wire [63:0]      spc908_rtl_pc;
    wire sas_m908;
    reg [63:0] spc908_phy_pc_w;

    

    reg spc909_inst_done;
    wire [1:0]   spc909_thread_id;
    wire [63:0]      spc909_rtl_pc;
    wire sas_m909;
    reg [63:0] spc909_phy_pc_w;

    

    reg spc910_inst_done;
    wire [1:0]   spc910_thread_id;
    wire [63:0]      spc910_rtl_pc;
    wire sas_m910;
    reg [63:0] spc910_phy_pc_w;

    

    reg spc911_inst_done;
    wire [1:0]   spc911_thread_id;
    wire [63:0]      spc911_rtl_pc;
    wire sas_m911;
    reg [63:0] spc911_phy_pc_w;

    

    reg spc912_inst_done;
    wire [1:0]   spc912_thread_id;
    wire [63:0]      spc912_rtl_pc;
    wire sas_m912;
    reg [63:0] spc912_phy_pc_w;

    

    reg spc913_inst_done;
    wire [1:0]   spc913_thread_id;
    wire [63:0]      spc913_rtl_pc;
    wire sas_m913;
    reg [63:0] spc913_phy_pc_w;

    

    reg spc914_inst_done;
    wire [1:0]   spc914_thread_id;
    wire [63:0]      spc914_rtl_pc;
    wire sas_m914;
    reg [63:0] spc914_phy_pc_w;

    

    reg spc915_inst_done;
    wire [1:0]   spc915_thread_id;
    wire [63:0]      spc915_rtl_pc;
    wire sas_m915;
    reg [63:0] spc915_phy_pc_w;

    

    reg spc916_inst_done;
    wire [1:0]   spc916_thread_id;
    wire [63:0]      spc916_rtl_pc;
    wire sas_m916;
    reg [63:0] spc916_phy_pc_w;

    

    reg spc917_inst_done;
    wire [1:0]   spc917_thread_id;
    wire [63:0]      spc917_rtl_pc;
    wire sas_m917;
    reg [63:0] spc917_phy_pc_w;

    

    reg spc918_inst_done;
    wire [1:0]   spc918_thread_id;
    wire [63:0]      spc918_rtl_pc;
    wire sas_m918;
    reg [63:0] spc918_phy_pc_w;

    

    reg spc919_inst_done;
    wire [1:0]   spc919_thread_id;
    wire [63:0]      spc919_rtl_pc;
    wire sas_m919;
    reg [63:0] spc919_phy_pc_w;

    

    reg spc920_inst_done;
    wire [1:0]   spc920_thread_id;
    wire [63:0]      spc920_rtl_pc;
    wire sas_m920;
    reg [63:0] spc920_phy_pc_w;

    

    reg spc921_inst_done;
    wire [1:0]   spc921_thread_id;
    wire [63:0]      spc921_rtl_pc;
    wire sas_m921;
    reg [63:0] spc921_phy_pc_w;

    

    reg spc922_inst_done;
    wire [1:0]   spc922_thread_id;
    wire [63:0]      spc922_rtl_pc;
    wire sas_m922;
    reg [63:0] spc922_phy_pc_w;

    

    reg spc923_inst_done;
    wire [1:0]   spc923_thread_id;
    wire [63:0]      spc923_rtl_pc;
    wire sas_m923;
    reg [63:0] spc923_phy_pc_w;

    

    reg spc924_inst_done;
    wire [1:0]   spc924_thread_id;
    wire [63:0]      spc924_rtl_pc;
    wire sas_m924;
    reg [63:0] spc924_phy_pc_w;

    

    reg spc925_inst_done;
    wire [1:0]   spc925_thread_id;
    wire [63:0]      spc925_rtl_pc;
    wire sas_m925;
    reg [63:0] spc925_phy_pc_w;

    

    reg spc926_inst_done;
    wire [1:0]   spc926_thread_id;
    wire [63:0]      spc926_rtl_pc;
    wire sas_m926;
    reg [63:0] spc926_phy_pc_w;

    

    reg spc927_inst_done;
    wire [1:0]   spc927_thread_id;
    wire [63:0]      spc927_rtl_pc;
    wire sas_m927;
    reg [63:0] spc927_phy_pc_w;

    

    reg spc928_inst_done;
    wire [1:0]   spc928_thread_id;
    wire [63:0]      spc928_rtl_pc;
    wire sas_m928;
    reg [63:0] spc928_phy_pc_w;

    

    reg spc929_inst_done;
    wire [1:0]   spc929_thread_id;
    wire [63:0]      spc929_rtl_pc;
    wire sas_m929;
    reg [63:0] spc929_phy_pc_w;

    

    reg spc930_inst_done;
    wire [1:0]   spc930_thread_id;
    wire [63:0]      spc930_rtl_pc;
    wire sas_m930;
    reg [63:0] spc930_phy_pc_w;

    

    reg spc931_inst_done;
    wire [1:0]   spc931_thread_id;
    wire [63:0]      spc931_rtl_pc;
    wire sas_m931;
    reg [63:0] spc931_phy_pc_w;

    

    reg spc932_inst_done;
    wire [1:0]   spc932_thread_id;
    wire [63:0]      spc932_rtl_pc;
    wire sas_m932;
    reg [63:0] spc932_phy_pc_w;

    

    reg spc933_inst_done;
    wire [1:0]   spc933_thread_id;
    wire [63:0]      spc933_rtl_pc;
    wire sas_m933;
    reg [63:0] spc933_phy_pc_w;

    

    reg spc934_inst_done;
    wire [1:0]   spc934_thread_id;
    wire [63:0]      spc934_rtl_pc;
    wire sas_m934;
    reg [63:0] spc934_phy_pc_w;

    

    reg spc935_inst_done;
    wire [1:0]   spc935_thread_id;
    wire [63:0]      spc935_rtl_pc;
    wire sas_m935;
    reg [63:0] spc935_phy_pc_w;

    

    reg spc936_inst_done;
    wire [1:0]   spc936_thread_id;
    wire [63:0]      spc936_rtl_pc;
    wire sas_m936;
    reg [63:0] spc936_phy_pc_w;

    

    reg spc937_inst_done;
    wire [1:0]   spc937_thread_id;
    wire [63:0]      spc937_rtl_pc;
    wire sas_m937;
    reg [63:0] spc937_phy_pc_w;

    

    reg spc938_inst_done;
    wire [1:0]   spc938_thread_id;
    wire [63:0]      spc938_rtl_pc;
    wire sas_m938;
    reg [63:0] spc938_phy_pc_w;

    

    reg spc939_inst_done;
    wire [1:0]   spc939_thread_id;
    wire [63:0]      spc939_rtl_pc;
    wire sas_m939;
    reg [63:0] spc939_phy_pc_w;

    

    reg spc940_inst_done;
    wire [1:0]   spc940_thread_id;
    wire [63:0]      spc940_rtl_pc;
    wire sas_m940;
    reg [63:0] spc940_phy_pc_w;

    

    reg spc941_inst_done;
    wire [1:0]   spc941_thread_id;
    wire [63:0]      spc941_rtl_pc;
    wire sas_m941;
    reg [63:0] spc941_phy_pc_w;

    

    reg spc942_inst_done;
    wire [1:0]   spc942_thread_id;
    wire [63:0]      spc942_rtl_pc;
    wire sas_m942;
    reg [63:0] spc942_phy_pc_w;

    

    reg spc943_inst_done;
    wire [1:0]   spc943_thread_id;
    wire [63:0]      spc943_rtl_pc;
    wire sas_m943;
    reg [63:0] spc943_phy_pc_w;

    

    reg spc944_inst_done;
    wire [1:0]   spc944_thread_id;
    wire [63:0]      spc944_rtl_pc;
    wire sas_m944;
    reg [63:0] spc944_phy_pc_w;

    

    reg spc945_inst_done;
    wire [1:0]   spc945_thread_id;
    wire [63:0]      spc945_rtl_pc;
    wire sas_m945;
    reg [63:0] spc945_phy_pc_w;

    

    reg spc946_inst_done;
    wire [1:0]   spc946_thread_id;
    wire [63:0]      spc946_rtl_pc;
    wire sas_m946;
    reg [63:0] spc946_phy_pc_w;

    

    reg spc947_inst_done;
    wire [1:0]   spc947_thread_id;
    wire [63:0]      spc947_rtl_pc;
    wire sas_m947;
    reg [63:0] spc947_phy_pc_w;

    

    reg spc948_inst_done;
    wire [1:0]   spc948_thread_id;
    wire [63:0]      spc948_rtl_pc;
    wire sas_m948;
    reg [63:0] spc948_phy_pc_w;

    

    reg spc949_inst_done;
    wire [1:0]   spc949_thread_id;
    wire [63:0]      spc949_rtl_pc;
    wire sas_m949;
    reg [63:0] spc949_phy_pc_w;

    

    reg spc950_inst_done;
    wire [1:0]   spc950_thread_id;
    wire [63:0]      spc950_rtl_pc;
    wire sas_m950;
    reg [63:0] spc950_phy_pc_w;

    

    reg spc951_inst_done;
    wire [1:0]   spc951_thread_id;
    wire [63:0]      spc951_rtl_pc;
    wire sas_m951;
    reg [63:0] spc951_phy_pc_w;

    

    reg spc952_inst_done;
    wire [1:0]   spc952_thread_id;
    wire [63:0]      spc952_rtl_pc;
    wire sas_m952;
    reg [63:0] spc952_phy_pc_w;

    

    reg spc953_inst_done;
    wire [1:0]   spc953_thread_id;
    wire [63:0]      spc953_rtl_pc;
    wire sas_m953;
    reg [63:0] spc953_phy_pc_w;

    

    reg spc954_inst_done;
    wire [1:0]   spc954_thread_id;
    wire [63:0]      spc954_rtl_pc;
    wire sas_m954;
    reg [63:0] spc954_phy_pc_w;

    

    reg spc955_inst_done;
    wire [1:0]   spc955_thread_id;
    wire [63:0]      spc955_rtl_pc;
    wire sas_m955;
    reg [63:0] spc955_phy_pc_w;

    

    reg spc956_inst_done;
    wire [1:0]   spc956_thread_id;
    wire [63:0]      spc956_rtl_pc;
    wire sas_m956;
    reg [63:0] spc956_phy_pc_w;

    

    reg spc957_inst_done;
    wire [1:0]   spc957_thread_id;
    wire [63:0]      spc957_rtl_pc;
    wire sas_m957;
    reg [63:0] spc957_phy_pc_w;

    

    reg spc958_inst_done;
    wire [1:0]   spc958_thread_id;
    wire [63:0]      spc958_rtl_pc;
    wire sas_m958;
    reg [63:0] spc958_phy_pc_w;

    

    reg spc959_inst_done;
    wire [1:0]   spc959_thread_id;
    wire [63:0]      spc959_rtl_pc;
    wire sas_m959;
    reg [63:0] spc959_phy_pc_w;

    

    reg spc960_inst_done;
    wire [1:0]   spc960_thread_id;
    wire [63:0]      spc960_rtl_pc;
    wire sas_m960;
    reg [63:0] spc960_phy_pc_w;

    

    reg spc961_inst_done;
    wire [1:0]   spc961_thread_id;
    wire [63:0]      spc961_rtl_pc;
    wire sas_m961;
    reg [63:0] spc961_phy_pc_w;

    

    reg spc962_inst_done;
    wire [1:0]   spc962_thread_id;
    wire [63:0]      spc962_rtl_pc;
    wire sas_m962;
    reg [63:0] spc962_phy_pc_w;

    

    reg spc963_inst_done;
    wire [1:0]   spc963_thread_id;
    wire [63:0]      spc963_rtl_pc;
    wire sas_m963;
    reg [63:0] spc963_phy_pc_w;

    

    reg spc964_inst_done;
    wire [1:0]   spc964_thread_id;
    wire [63:0]      spc964_rtl_pc;
    wire sas_m964;
    reg [63:0] spc964_phy_pc_w;

    

    reg spc965_inst_done;
    wire [1:0]   spc965_thread_id;
    wire [63:0]      spc965_rtl_pc;
    wire sas_m965;
    reg [63:0] spc965_phy_pc_w;

    

    reg spc966_inst_done;
    wire [1:0]   spc966_thread_id;
    wire [63:0]      spc966_rtl_pc;
    wire sas_m966;
    reg [63:0] spc966_phy_pc_w;

    

    reg spc967_inst_done;
    wire [1:0]   spc967_thread_id;
    wire [63:0]      spc967_rtl_pc;
    wire sas_m967;
    reg [63:0] spc967_phy_pc_w;

    

    reg spc968_inst_done;
    wire [1:0]   spc968_thread_id;
    wire [63:0]      spc968_rtl_pc;
    wire sas_m968;
    reg [63:0] spc968_phy_pc_w;

    

    reg spc969_inst_done;
    wire [1:0]   spc969_thread_id;
    wire [63:0]      spc969_rtl_pc;
    wire sas_m969;
    reg [63:0] spc969_phy_pc_w;

    

    reg spc970_inst_done;
    wire [1:0]   spc970_thread_id;
    wire [63:0]      spc970_rtl_pc;
    wire sas_m970;
    reg [63:0] spc970_phy_pc_w;

    

    reg spc971_inst_done;
    wire [1:0]   spc971_thread_id;
    wire [63:0]      spc971_rtl_pc;
    wire sas_m971;
    reg [63:0] spc971_phy_pc_w;

    

    reg spc972_inst_done;
    wire [1:0]   spc972_thread_id;
    wire [63:0]      spc972_rtl_pc;
    wire sas_m972;
    reg [63:0] spc972_phy_pc_w;

    

    reg spc973_inst_done;
    wire [1:0]   spc973_thread_id;
    wire [63:0]      spc973_rtl_pc;
    wire sas_m973;
    reg [63:0] spc973_phy_pc_w;

    

    reg spc974_inst_done;
    wire [1:0]   spc974_thread_id;
    wire [63:0]      spc974_rtl_pc;
    wire sas_m974;
    reg [63:0] spc974_phy_pc_w;

    

    reg spc975_inst_done;
    wire [1:0]   spc975_thread_id;
    wire [63:0]      spc975_rtl_pc;
    wire sas_m975;
    reg [63:0] spc975_phy_pc_w;

    

    reg spc976_inst_done;
    wire [1:0]   spc976_thread_id;
    wire [63:0]      spc976_rtl_pc;
    wire sas_m976;
    reg [63:0] spc976_phy_pc_w;

    

    reg spc977_inst_done;
    wire [1:0]   spc977_thread_id;
    wire [63:0]      spc977_rtl_pc;
    wire sas_m977;
    reg [63:0] spc977_phy_pc_w;

    

    reg spc978_inst_done;
    wire [1:0]   spc978_thread_id;
    wire [63:0]      spc978_rtl_pc;
    wire sas_m978;
    reg [63:0] spc978_phy_pc_w;

    

    reg spc979_inst_done;
    wire [1:0]   spc979_thread_id;
    wire [63:0]      spc979_rtl_pc;
    wire sas_m979;
    reg [63:0] spc979_phy_pc_w;

    

    reg spc980_inst_done;
    wire [1:0]   spc980_thread_id;
    wire [63:0]      spc980_rtl_pc;
    wire sas_m980;
    reg [63:0] spc980_phy_pc_w;

    

    reg spc981_inst_done;
    wire [1:0]   spc981_thread_id;
    wire [63:0]      spc981_rtl_pc;
    wire sas_m981;
    reg [63:0] spc981_phy_pc_w;

    

    reg spc982_inst_done;
    wire [1:0]   spc982_thread_id;
    wire [63:0]      spc982_rtl_pc;
    wire sas_m982;
    reg [63:0] spc982_phy_pc_w;

    

    reg spc983_inst_done;
    wire [1:0]   spc983_thread_id;
    wire [63:0]      spc983_rtl_pc;
    wire sas_m983;
    reg [63:0] spc983_phy_pc_w;

    

    reg spc984_inst_done;
    wire [1:0]   spc984_thread_id;
    wire [63:0]      spc984_rtl_pc;
    wire sas_m984;
    reg [63:0] spc984_phy_pc_w;

    

    reg spc985_inst_done;
    wire [1:0]   spc985_thread_id;
    wire [63:0]      spc985_rtl_pc;
    wire sas_m985;
    reg [63:0] spc985_phy_pc_w;

    

    reg spc986_inst_done;
    wire [1:0]   spc986_thread_id;
    wire [63:0]      spc986_rtl_pc;
    wire sas_m986;
    reg [63:0] spc986_phy_pc_w;

    

    reg spc987_inst_done;
    wire [1:0]   spc987_thread_id;
    wire [63:0]      spc987_rtl_pc;
    wire sas_m987;
    reg [63:0] spc987_phy_pc_w;

    

    reg spc988_inst_done;
    wire [1:0]   spc988_thread_id;
    wire [63:0]      spc988_rtl_pc;
    wire sas_m988;
    reg [63:0] spc988_phy_pc_w;

    

    reg spc989_inst_done;
    wire [1:0]   spc989_thread_id;
    wire [63:0]      spc989_rtl_pc;
    wire sas_m989;
    reg [63:0] spc989_phy_pc_w;

    

    reg spc990_inst_done;
    wire [1:0]   spc990_thread_id;
    wire [63:0]      spc990_rtl_pc;
    wire sas_m990;
    reg [63:0] spc990_phy_pc_w;

    

    reg spc991_inst_done;
    wire [1:0]   spc991_thread_id;
    wire [63:0]      spc991_rtl_pc;
    wire sas_m991;
    reg [63:0] spc991_phy_pc_w;

    

    reg spc992_inst_done;
    wire [1:0]   spc992_thread_id;
    wire [63:0]      spc992_rtl_pc;
    wire sas_m992;
    reg [63:0] spc992_phy_pc_w;

    

    reg spc993_inst_done;
    wire [1:0]   spc993_thread_id;
    wire [63:0]      spc993_rtl_pc;
    wire sas_m993;
    reg [63:0] spc993_phy_pc_w;

    

    reg spc994_inst_done;
    wire [1:0]   spc994_thread_id;
    wire [63:0]      spc994_rtl_pc;
    wire sas_m994;
    reg [63:0] spc994_phy_pc_w;

    

    reg spc995_inst_done;
    wire [1:0]   spc995_thread_id;
    wire [63:0]      spc995_rtl_pc;
    wire sas_m995;
    reg [63:0] spc995_phy_pc_w;

    

    reg spc996_inst_done;
    wire [1:0]   spc996_thread_id;
    wire [63:0]      spc996_rtl_pc;
    wire sas_m996;
    reg [63:0] spc996_phy_pc_w;

    

    reg spc997_inst_done;
    wire [1:0]   spc997_thread_id;
    wire [63:0]      spc997_rtl_pc;
    wire sas_m997;
    reg [63:0] spc997_phy_pc_w;

    

    reg spc998_inst_done;
    wire [1:0]   spc998_thread_id;
    wire [63:0]      spc998_rtl_pc;
    wire sas_m998;
    reg [63:0] spc998_phy_pc_w;

    

    reg spc999_inst_done;
    wire [1:0]   spc999_thread_id;
    wire [63:0]      spc999_rtl_pc;
    wire sas_m999;
    reg [63:0] spc999_phy_pc_w;

    

    reg spc1000_inst_done;
    wire [1:0]   spc1000_thread_id;
    wire [63:0]      spc1000_rtl_pc;
    wire sas_m1000;
    reg [63:0] spc1000_phy_pc_w;

    

    reg spc1001_inst_done;
    wire [1:0]   spc1001_thread_id;
    wire [63:0]      spc1001_rtl_pc;
    wire sas_m1001;
    reg [63:0] spc1001_phy_pc_w;

    

    reg spc1002_inst_done;
    wire [1:0]   spc1002_thread_id;
    wire [63:0]      spc1002_rtl_pc;
    wire sas_m1002;
    reg [63:0] spc1002_phy_pc_w;

    

    reg spc1003_inst_done;
    wire [1:0]   spc1003_thread_id;
    wire [63:0]      spc1003_rtl_pc;
    wire sas_m1003;
    reg [63:0] spc1003_phy_pc_w;

    

    reg spc1004_inst_done;
    wire [1:0]   spc1004_thread_id;
    wire [63:0]      spc1004_rtl_pc;
    wire sas_m1004;
    reg [63:0] spc1004_phy_pc_w;

    

    reg spc1005_inst_done;
    wire [1:0]   spc1005_thread_id;
    wire [63:0]      spc1005_rtl_pc;
    wire sas_m1005;
    reg [63:0] spc1005_phy_pc_w;

    

    reg spc1006_inst_done;
    wire [1:0]   spc1006_thread_id;
    wire [63:0]      spc1006_rtl_pc;
    wire sas_m1006;
    reg [63:0] spc1006_phy_pc_w;

    

    reg spc1007_inst_done;
    wire [1:0]   spc1007_thread_id;
    wire [63:0]      spc1007_rtl_pc;
    wire sas_m1007;
    reg [63:0] spc1007_phy_pc_w;

    

    reg spc1008_inst_done;
    wire [1:0]   spc1008_thread_id;
    wire [63:0]      spc1008_rtl_pc;
    wire sas_m1008;
    reg [63:0] spc1008_phy_pc_w;

    

    reg spc1009_inst_done;
    wire [1:0]   spc1009_thread_id;
    wire [63:0]      spc1009_rtl_pc;
    wire sas_m1009;
    reg [63:0] spc1009_phy_pc_w;

    

    reg spc1010_inst_done;
    wire [1:0]   spc1010_thread_id;
    wire [63:0]      spc1010_rtl_pc;
    wire sas_m1010;
    reg [63:0] spc1010_phy_pc_w;

    

    reg spc1011_inst_done;
    wire [1:0]   spc1011_thread_id;
    wire [63:0]      spc1011_rtl_pc;
    wire sas_m1011;
    reg [63:0] spc1011_phy_pc_w;

    

    reg spc1012_inst_done;
    wire [1:0]   spc1012_thread_id;
    wire [63:0]      spc1012_rtl_pc;
    wire sas_m1012;
    reg [63:0] spc1012_phy_pc_w;

    

    reg spc1013_inst_done;
    wire [1:0]   spc1013_thread_id;
    wire [63:0]      spc1013_rtl_pc;
    wire sas_m1013;
    reg [63:0] spc1013_phy_pc_w;

    

    reg spc1014_inst_done;
    wire [1:0]   spc1014_thread_id;
    wire [63:0]      spc1014_rtl_pc;
    wire sas_m1014;
    reg [63:0] spc1014_phy_pc_w;

    

    reg spc1015_inst_done;
    wire [1:0]   spc1015_thread_id;
    wire [63:0]      spc1015_rtl_pc;
    wire sas_m1015;
    reg [63:0] spc1015_phy_pc_w;

    

    reg spc1016_inst_done;
    wire [1:0]   spc1016_thread_id;
    wire [63:0]      spc1016_rtl_pc;
    wire sas_m1016;
    reg [63:0] spc1016_phy_pc_w;

    

    reg spc1017_inst_done;
    wire [1:0]   spc1017_thread_id;
    wire [63:0]      spc1017_rtl_pc;
    wire sas_m1017;
    reg [63:0] spc1017_phy_pc_w;

    

    reg spc1018_inst_done;
    wire [1:0]   spc1018_thread_id;
    wire [63:0]      spc1018_rtl_pc;
    wire sas_m1018;
    reg [63:0] spc1018_phy_pc_w;

    

    reg spc1019_inst_done;
    wire [1:0]   spc1019_thread_id;
    wire [63:0]      spc1019_rtl_pc;
    wire sas_m1019;
    reg [63:0] spc1019_phy_pc_w;

    

    reg spc1020_inst_done;
    wire [1:0]   spc1020_thread_id;
    wire [63:0]      spc1020_rtl_pc;
    wire sas_m1020;
    reg [63:0] spc1020_phy_pc_w;

    

    reg spc1021_inst_done;
    wire [1:0]   spc1021_thread_id;
    wire [63:0]      spc1021_rtl_pc;
    wire sas_m1021;
    reg [63:0] spc1021_phy_pc_w;

    

    reg spc1022_inst_done;
    wire [1:0]   spc1022_thread_id;
    wire [63:0]      spc1022_rtl_pc;
    wire sas_m1022;
    reg [63:0] spc1022_phy_pc_w;

    

    reg spc1023_inst_done;
    wire [1:0]   spc1023_thread_id;
    wire [63:0]      spc1023_rtl_pc;
    wire sas_m1023;
    reg [63:0] spc1023_phy_pc_w;

    


integer      good_trap_count;
integer      bad_trap_count;
reg         local_diag_done;

//use this for the second reset.
initial begin
    local_diag_done = 0;

    good_trap_exists = {`GOOD_TRAP_COUNTER{1'b0}};
    bad_trap_exists = {`GOOD_TRAP_COUNTER{1'b0}};
end
//-----------------------------------------------------------

`ifdef INCLUDE_SAS_TASKS
task get_thread_status;
    begin
    thread_status[0] = `IFUPATH0.swl.thr0_state;
thread_status[1] = `IFUPATH0.swl.thr1_state;
thread_status[2] = `IFUPATH0.swl.thr2_state;
thread_status[3] = `IFUPATH0.swl.thr3_state;
thread_status[4] = `IFUPATH1.swl.thr0_state;
thread_status[5] = `IFUPATH1.swl.thr1_state;
thread_status[6] = `IFUPATH1.swl.thr2_state;
thread_status[7] = `IFUPATH1.swl.thr3_state;
thread_status[8] = `IFUPATH2.swl.thr0_state;
thread_status[9] = `IFUPATH2.swl.thr1_state;
thread_status[10] = `IFUPATH2.swl.thr2_state;
thread_status[11] = `IFUPATH2.swl.thr3_state;
thread_status[12] = `IFUPATH3.swl.thr0_state;
thread_status[13] = `IFUPATH3.swl.thr1_state;
thread_status[14] = `IFUPATH3.swl.thr2_state;
thread_status[15] = `IFUPATH3.swl.thr3_state;
thread_status[16] = `IFUPATH4.swl.thr0_state;
thread_status[17] = `IFUPATH4.swl.thr1_state;
thread_status[18] = `IFUPATH4.swl.thr2_state;
thread_status[19] = `IFUPATH4.swl.thr3_state;
thread_status[20] = `IFUPATH5.swl.thr0_state;
thread_status[21] = `IFUPATH5.swl.thr1_state;
thread_status[22] = `IFUPATH5.swl.thr2_state;
thread_status[23] = `IFUPATH5.swl.thr3_state;
thread_status[24] = `IFUPATH6.swl.thr0_state;
thread_status[25] = `IFUPATH6.swl.thr1_state;
thread_status[26] = `IFUPATH6.swl.thr2_state;
thread_status[27] = `IFUPATH6.swl.thr3_state;
thread_status[28] = `IFUPATH7.swl.thr0_state;
thread_status[29] = `IFUPATH7.swl.thr1_state;
thread_status[30] = `IFUPATH7.swl.thr2_state;
thread_status[31] = `IFUPATH7.swl.thr3_state;
thread_status[32] = `IFUPATH8.swl.thr0_state;
thread_status[33] = `IFUPATH8.swl.thr1_state;
thread_status[34] = `IFUPATH8.swl.thr2_state;
thread_status[35] = `IFUPATH8.swl.thr3_state;
thread_status[36] = `IFUPATH9.swl.thr0_state;
thread_status[37] = `IFUPATH9.swl.thr1_state;
thread_status[38] = `IFUPATH9.swl.thr2_state;
thread_status[39] = `IFUPATH9.swl.thr3_state;
thread_status[40] = `IFUPATH10.swl.thr0_state;
thread_status[41] = `IFUPATH10.swl.thr1_state;
thread_status[42] = `IFUPATH10.swl.thr2_state;
thread_status[43] = `IFUPATH10.swl.thr3_state;
thread_status[44] = `IFUPATH11.swl.thr0_state;
thread_status[45] = `IFUPATH11.swl.thr1_state;
thread_status[46] = `IFUPATH11.swl.thr2_state;
thread_status[47] = `IFUPATH11.swl.thr3_state;
thread_status[48] = `IFUPATH12.swl.thr0_state;
thread_status[49] = `IFUPATH12.swl.thr1_state;
thread_status[50] = `IFUPATH12.swl.thr2_state;
thread_status[51] = `IFUPATH12.swl.thr3_state;
thread_status[52] = `IFUPATH13.swl.thr0_state;
thread_status[53] = `IFUPATH13.swl.thr1_state;
thread_status[54] = `IFUPATH13.swl.thr2_state;
thread_status[55] = `IFUPATH13.swl.thr3_state;
thread_status[56] = `IFUPATH14.swl.thr0_state;
thread_status[57] = `IFUPATH14.swl.thr1_state;
thread_status[58] = `IFUPATH14.swl.thr2_state;
thread_status[59] = `IFUPATH14.swl.thr3_state;
thread_status[60] = `IFUPATH15.swl.thr0_state;
thread_status[61] = `IFUPATH15.swl.thr1_state;
thread_status[62] = `IFUPATH15.swl.thr2_state;
thread_status[63] = `IFUPATH15.swl.thr3_state;
thread_status[64] = `IFUPATH16.swl.thr0_state;
thread_status[65] = `IFUPATH16.swl.thr1_state;
thread_status[66] = `IFUPATH16.swl.thr2_state;
thread_status[67] = `IFUPATH16.swl.thr3_state;
thread_status[68] = `IFUPATH17.swl.thr0_state;
thread_status[69] = `IFUPATH17.swl.thr1_state;
thread_status[70] = `IFUPATH17.swl.thr2_state;
thread_status[71] = `IFUPATH17.swl.thr3_state;
thread_status[72] = `IFUPATH18.swl.thr0_state;
thread_status[73] = `IFUPATH18.swl.thr1_state;
thread_status[74] = `IFUPATH18.swl.thr2_state;
thread_status[75] = `IFUPATH18.swl.thr3_state;
thread_status[76] = `IFUPATH19.swl.thr0_state;
thread_status[77] = `IFUPATH19.swl.thr1_state;
thread_status[78] = `IFUPATH19.swl.thr2_state;
thread_status[79] = `IFUPATH19.swl.thr3_state;
thread_status[80] = `IFUPATH20.swl.thr0_state;
thread_status[81] = `IFUPATH20.swl.thr1_state;
thread_status[82] = `IFUPATH20.swl.thr2_state;
thread_status[83] = `IFUPATH20.swl.thr3_state;
thread_status[84] = `IFUPATH21.swl.thr0_state;
thread_status[85] = `IFUPATH21.swl.thr1_state;
thread_status[86] = `IFUPATH21.swl.thr2_state;
thread_status[87] = `IFUPATH21.swl.thr3_state;
thread_status[88] = `IFUPATH22.swl.thr0_state;
thread_status[89] = `IFUPATH22.swl.thr1_state;
thread_status[90] = `IFUPATH22.swl.thr2_state;
thread_status[91] = `IFUPATH22.swl.thr3_state;
thread_status[92] = `IFUPATH23.swl.thr0_state;
thread_status[93] = `IFUPATH23.swl.thr1_state;
thread_status[94] = `IFUPATH23.swl.thr2_state;
thread_status[95] = `IFUPATH23.swl.thr3_state;
thread_status[96] = `IFUPATH24.swl.thr0_state;
thread_status[97] = `IFUPATH24.swl.thr1_state;
thread_status[98] = `IFUPATH24.swl.thr2_state;
thread_status[99] = `IFUPATH24.swl.thr3_state;
thread_status[100] = `IFUPATH25.swl.thr0_state;
thread_status[101] = `IFUPATH25.swl.thr1_state;
thread_status[102] = `IFUPATH25.swl.thr2_state;
thread_status[103] = `IFUPATH25.swl.thr3_state;
thread_status[104] = `IFUPATH26.swl.thr0_state;
thread_status[105] = `IFUPATH26.swl.thr1_state;
thread_status[106] = `IFUPATH26.swl.thr2_state;
thread_status[107] = `IFUPATH26.swl.thr3_state;
thread_status[108] = `IFUPATH27.swl.thr0_state;
thread_status[109] = `IFUPATH27.swl.thr1_state;
thread_status[110] = `IFUPATH27.swl.thr2_state;
thread_status[111] = `IFUPATH27.swl.thr3_state;
thread_status[112] = `IFUPATH28.swl.thr0_state;
thread_status[113] = `IFUPATH28.swl.thr1_state;
thread_status[114] = `IFUPATH28.swl.thr2_state;
thread_status[115] = `IFUPATH28.swl.thr3_state;
thread_status[116] = `IFUPATH29.swl.thr0_state;
thread_status[117] = `IFUPATH29.swl.thr1_state;
thread_status[118] = `IFUPATH29.swl.thr2_state;
thread_status[119] = `IFUPATH29.swl.thr3_state;
thread_status[120] = `IFUPATH30.swl.thr0_state;
thread_status[121] = `IFUPATH30.swl.thr1_state;
thread_status[122] = `IFUPATH30.swl.thr2_state;
thread_status[123] = `IFUPATH30.swl.thr3_state;
thread_status[124] = `IFUPATH31.swl.thr0_state;
thread_status[125] = `IFUPATH31.swl.thr1_state;
thread_status[126] = `IFUPATH31.swl.thr2_state;
thread_status[127] = `IFUPATH31.swl.thr3_state;
thread_status[128] = `IFUPATH32.swl.thr0_state;
thread_status[129] = `IFUPATH32.swl.thr1_state;
thread_status[130] = `IFUPATH32.swl.thr2_state;
thread_status[131] = `IFUPATH32.swl.thr3_state;
thread_status[132] = `IFUPATH33.swl.thr0_state;
thread_status[133] = `IFUPATH33.swl.thr1_state;
thread_status[134] = `IFUPATH33.swl.thr2_state;
thread_status[135] = `IFUPATH33.swl.thr3_state;
thread_status[136] = `IFUPATH34.swl.thr0_state;
thread_status[137] = `IFUPATH34.swl.thr1_state;
thread_status[138] = `IFUPATH34.swl.thr2_state;
thread_status[139] = `IFUPATH34.swl.thr3_state;
thread_status[140] = `IFUPATH35.swl.thr0_state;
thread_status[141] = `IFUPATH35.swl.thr1_state;
thread_status[142] = `IFUPATH35.swl.thr2_state;
thread_status[143] = `IFUPATH35.swl.thr3_state;
thread_status[144] = `IFUPATH36.swl.thr0_state;
thread_status[145] = `IFUPATH36.swl.thr1_state;
thread_status[146] = `IFUPATH36.swl.thr2_state;
thread_status[147] = `IFUPATH36.swl.thr3_state;
thread_status[148] = `IFUPATH37.swl.thr0_state;
thread_status[149] = `IFUPATH37.swl.thr1_state;
thread_status[150] = `IFUPATH37.swl.thr2_state;
thread_status[151] = `IFUPATH37.swl.thr3_state;
thread_status[152] = `IFUPATH38.swl.thr0_state;
thread_status[153] = `IFUPATH38.swl.thr1_state;
thread_status[154] = `IFUPATH38.swl.thr2_state;
thread_status[155] = `IFUPATH38.swl.thr3_state;
thread_status[156] = `IFUPATH39.swl.thr0_state;
thread_status[157] = `IFUPATH39.swl.thr1_state;
thread_status[158] = `IFUPATH39.swl.thr2_state;
thread_status[159] = `IFUPATH39.swl.thr3_state;
thread_status[160] = `IFUPATH40.swl.thr0_state;
thread_status[161] = `IFUPATH40.swl.thr1_state;
thread_status[162] = `IFUPATH40.swl.thr2_state;
thread_status[163] = `IFUPATH40.swl.thr3_state;
thread_status[164] = `IFUPATH41.swl.thr0_state;
thread_status[165] = `IFUPATH41.swl.thr1_state;
thread_status[166] = `IFUPATH41.swl.thr2_state;
thread_status[167] = `IFUPATH41.swl.thr3_state;
thread_status[168] = `IFUPATH42.swl.thr0_state;
thread_status[169] = `IFUPATH42.swl.thr1_state;
thread_status[170] = `IFUPATH42.swl.thr2_state;
thread_status[171] = `IFUPATH42.swl.thr3_state;
thread_status[172] = `IFUPATH43.swl.thr0_state;
thread_status[173] = `IFUPATH43.swl.thr1_state;
thread_status[174] = `IFUPATH43.swl.thr2_state;
thread_status[175] = `IFUPATH43.swl.thr3_state;
thread_status[176] = `IFUPATH44.swl.thr0_state;
thread_status[177] = `IFUPATH44.swl.thr1_state;
thread_status[178] = `IFUPATH44.swl.thr2_state;
thread_status[179] = `IFUPATH44.swl.thr3_state;
thread_status[180] = `IFUPATH45.swl.thr0_state;
thread_status[181] = `IFUPATH45.swl.thr1_state;
thread_status[182] = `IFUPATH45.swl.thr2_state;
thread_status[183] = `IFUPATH45.swl.thr3_state;
thread_status[184] = `IFUPATH46.swl.thr0_state;
thread_status[185] = `IFUPATH46.swl.thr1_state;
thread_status[186] = `IFUPATH46.swl.thr2_state;
thread_status[187] = `IFUPATH46.swl.thr3_state;
thread_status[188] = `IFUPATH47.swl.thr0_state;
thread_status[189] = `IFUPATH47.swl.thr1_state;
thread_status[190] = `IFUPATH47.swl.thr2_state;
thread_status[191] = `IFUPATH47.swl.thr3_state;
thread_status[192] = `IFUPATH48.swl.thr0_state;
thread_status[193] = `IFUPATH48.swl.thr1_state;
thread_status[194] = `IFUPATH48.swl.thr2_state;
thread_status[195] = `IFUPATH48.swl.thr3_state;
thread_status[196] = `IFUPATH49.swl.thr0_state;
thread_status[197] = `IFUPATH49.swl.thr1_state;
thread_status[198] = `IFUPATH49.swl.thr2_state;
thread_status[199] = `IFUPATH49.swl.thr3_state;
thread_status[200] = `IFUPATH50.swl.thr0_state;
thread_status[201] = `IFUPATH50.swl.thr1_state;
thread_status[202] = `IFUPATH50.swl.thr2_state;
thread_status[203] = `IFUPATH50.swl.thr3_state;
thread_status[204] = `IFUPATH51.swl.thr0_state;
thread_status[205] = `IFUPATH51.swl.thr1_state;
thread_status[206] = `IFUPATH51.swl.thr2_state;
thread_status[207] = `IFUPATH51.swl.thr3_state;
thread_status[208] = `IFUPATH52.swl.thr0_state;
thread_status[209] = `IFUPATH52.swl.thr1_state;
thread_status[210] = `IFUPATH52.swl.thr2_state;
thread_status[211] = `IFUPATH52.swl.thr3_state;
thread_status[212] = `IFUPATH53.swl.thr0_state;
thread_status[213] = `IFUPATH53.swl.thr1_state;
thread_status[214] = `IFUPATH53.swl.thr2_state;
thread_status[215] = `IFUPATH53.swl.thr3_state;
thread_status[216] = `IFUPATH54.swl.thr0_state;
thread_status[217] = `IFUPATH54.swl.thr1_state;
thread_status[218] = `IFUPATH54.swl.thr2_state;
thread_status[219] = `IFUPATH54.swl.thr3_state;
thread_status[220] = `IFUPATH55.swl.thr0_state;
thread_status[221] = `IFUPATH55.swl.thr1_state;
thread_status[222] = `IFUPATH55.swl.thr2_state;
thread_status[223] = `IFUPATH55.swl.thr3_state;
thread_status[224] = `IFUPATH56.swl.thr0_state;
thread_status[225] = `IFUPATH56.swl.thr1_state;
thread_status[226] = `IFUPATH56.swl.thr2_state;
thread_status[227] = `IFUPATH56.swl.thr3_state;
thread_status[228] = `IFUPATH57.swl.thr0_state;
thread_status[229] = `IFUPATH57.swl.thr1_state;
thread_status[230] = `IFUPATH57.swl.thr2_state;
thread_status[231] = `IFUPATH57.swl.thr3_state;
thread_status[232] = `IFUPATH58.swl.thr0_state;
thread_status[233] = `IFUPATH58.swl.thr1_state;
thread_status[234] = `IFUPATH58.swl.thr2_state;
thread_status[235] = `IFUPATH58.swl.thr3_state;
thread_status[236] = `IFUPATH59.swl.thr0_state;
thread_status[237] = `IFUPATH59.swl.thr1_state;
thread_status[238] = `IFUPATH59.swl.thr2_state;
thread_status[239] = `IFUPATH59.swl.thr3_state;
thread_status[240] = `IFUPATH60.swl.thr0_state;
thread_status[241] = `IFUPATH60.swl.thr1_state;
thread_status[242] = `IFUPATH60.swl.thr2_state;
thread_status[243] = `IFUPATH60.swl.thr3_state;
thread_status[244] = `IFUPATH61.swl.thr0_state;
thread_status[245] = `IFUPATH61.swl.thr1_state;
thread_status[246] = `IFUPATH61.swl.thr2_state;
thread_status[247] = `IFUPATH61.swl.thr3_state;
thread_status[248] = `IFUPATH62.swl.thr0_state;
thread_status[249] = `IFUPATH62.swl.thr1_state;
thread_status[250] = `IFUPATH62.swl.thr2_state;
thread_status[251] = `IFUPATH62.swl.thr3_state;
thread_status[252] = `IFUPATH63.swl.thr0_state;
thread_status[253] = `IFUPATH63.swl.thr1_state;
thread_status[254] = `IFUPATH63.swl.thr2_state;
thread_status[255] = `IFUPATH63.swl.thr3_state;
thread_status[256] = `IFUPATH64.swl.thr0_state;
thread_status[257] = `IFUPATH64.swl.thr1_state;
thread_status[258] = `IFUPATH64.swl.thr2_state;
thread_status[259] = `IFUPATH64.swl.thr3_state;
thread_status[260] = `IFUPATH65.swl.thr0_state;
thread_status[261] = `IFUPATH65.swl.thr1_state;
thread_status[262] = `IFUPATH65.swl.thr2_state;
thread_status[263] = `IFUPATH65.swl.thr3_state;
thread_status[264] = `IFUPATH66.swl.thr0_state;
thread_status[265] = `IFUPATH66.swl.thr1_state;
thread_status[266] = `IFUPATH66.swl.thr2_state;
thread_status[267] = `IFUPATH66.swl.thr3_state;
thread_status[268] = `IFUPATH67.swl.thr0_state;
thread_status[269] = `IFUPATH67.swl.thr1_state;
thread_status[270] = `IFUPATH67.swl.thr2_state;
thread_status[271] = `IFUPATH67.swl.thr3_state;
thread_status[272] = `IFUPATH68.swl.thr0_state;
thread_status[273] = `IFUPATH68.swl.thr1_state;
thread_status[274] = `IFUPATH68.swl.thr2_state;
thread_status[275] = `IFUPATH68.swl.thr3_state;
thread_status[276] = `IFUPATH69.swl.thr0_state;
thread_status[277] = `IFUPATH69.swl.thr1_state;
thread_status[278] = `IFUPATH69.swl.thr2_state;
thread_status[279] = `IFUPATH69.swl.thr3_state;
thread_status[280] = `IFUPATH70.swl.thr0_state;
thread_status[281] = `IFUPATH70.swl.thr1_state;
thread_status[282] = `IFUPATH70.swl.thr2_state;
thread_status[283] = `IFUPATH70.swl.thr3_state;
thread_status[284] = `IFUPATH71.swl.thr0_state;
thread_status[285] = `IFUPATH71.swl.thr1_state;
thread_status[286] = `IFUPATH71.swl.thr2_state;
thread_status[287] = `IFUPATH71.swl.thr3_state;
thread_status[288] = `IFUPATH72.swl.thr0_state;
thread_status[289] = `IFUPATH72.swl.thr1_state;
thread_status[290] = `IFUPATH72.swl.thr2_state;
thread_status[291] = `IFUPATH72.swl.thr3_state;
thread_status[292] = `IFUPATH73.swl.thr0_state;
thread_status[293] = `IFUPATH73.swl.thr1_state;
thread_status[294] = `IFUPATH73.swl.thr2_state;
thread_status[295] = `IFUPATH73.swl.thr3_state;
thread_status[296] = `IFUPATH74.swl.thr0_state;
thread_status[297] = `IFUPATH74.swl.thr1_state;
thread_status[298] = `IFUPATH74.swl.thr2_state;
thread_status[299] = `IFUPATH74.swl.thr3_state;
thread_status[300] = `IFUPATH75.swl.thr0_state;
thread_status[301] = `IFUPATH75.swl.thr1_state;
thread_status[302] = `IFUPATH75.swl.thr2_state;
thread_status[303] = `IFUPATH75.swl.thr3_state;
thread_status[304] = `IFUPATH76.swl.thr0_state;
thread_status[305] = `IFUPATH76.swl.thr1_state;
thread_status[306] = `IFUPATH76.swl.thr2_state;
thread_status[307] = `IFUPATH76.swl.thr3_state;
thread_status[308] = `IFUPATH77.swl.thr0_state;
thread_status[309] = `IFUPATH77.swl.thr1_state;
thread_status[310] = `IFUPATH77.swl.thr2_state;
thread_status[311] = `IFUPATH77.swl.thr3_state;
thread_status[312] = `IFUPATH78.swl.thr0_state;
thread_status[313] = `IFUPATH78.swl.thr1_state;
thread_status[314] = `IFUPATH78.swl.thr2_state;
thread_status[315] = `IFUPATH78.swl.thr3_state;
thread_status[316] = `IFUPATH79.swl.thr0_state;
thread_status[317] = `IFUPATH79.swl.thr1_state;
thread_status[318] = `IFUPATH79.swl.thr2_state;
thread_status[319] = `IFUPATH79.swl.thr3_state;
thread_status[320] = `IFUPATH80.swl.thr0_state;
thread_status[321] = `IFUPATH80.swl.thr1_state;
thread_status[322] = `IFUPATH80.swl.thr2_state;
thread_status[323] = `IFUPATH80.swl.thr3_state;
thread_status[324] = `IFUPATH81.swl.thr0_state;
thread_status[325] = `IFUPATH81.swl.thr1_state;
thread_status[326] = `IFUPATH81.swl.thr2_state;
thread_status[327] = `IFUPATH81.swl.thr3_state;
thread_status[328] = `IFUPATH82.swl.thr0_state;
thread_status[329] = `IFUPATH82.swl.thr1_state;
thread_status[330] = `IFUPATH82.swl.thr2_state;
thread_status[331] = `IFUPATH82.swl.thr3_state;
thread_status[332] = `IFUPATH83.swl.thr0_state;
thread_status[333] = `IFUPATH83.swl.thr1_state;
thread_status[334] = `IFUPATH83.swl.thr2_state;
thread_status[335] = `IFUPATH83.swl.thr3_state;
thread_status[336] = `IFUPATH84.swl.thr0_state;
thread_status[337] = `IFUPATH84.swl.thr1_state;
thread_status[338] = `IFUPATH84.swl.thr2_state;
thread_status[339] = `IFUPATH84.swl.thr3_state;
thread_status[340] = `IFUPATH85.swl.thr0_state;
thread_status[341] = `IFUPATH85.swl.thr1_state;
thread_status[342] = `IFUPATH85.swl.thr2_state;
thread_status[343] = `IFUPATH85.swl.thr3_state;
thread_status[344] = `IFUPATH86.swl.thr0_state;
thread_status[345] = `IFUPATH86.swl.thr1_state;
thread_status[346] = `IFUPATH86.swl.thr2_state;
thread_status[347] = `IFUPATH86.swl.thr3_state;
thread_status[348] = `IFUPATH87.swl.thr0_state;
thread_status[349] = `IFUPATH87.swl.thr1_state;
thread_status[350] = `IFUPATH87.swl.thr2_state;
thread_status[351] = `IFUPATH87.swl.thr3_state;
thread_status[352] = `IFUPATH88.swl.thr0_state;
thread_status[353] = `IFUPATH88.swl.thr1_state;
thread_status[354] = `IFUPATH88.swl.thr2_state;
thread_status[355] = `IFUPATH88.swl.thr3_state;
thread_status[356] = `IFUPATH89.swl.thr0_state;
thread_status[357] = `IFUPATH89.swl.thr1_state;
thread_status[358] = `IFUPATH89.swl.thr2_state;
thread_status[359] = `IFUPATH89.swl.thr3_state;
thread_status[360] = `IFUPATH90.swl.thr0_state;
thread_status[361] = `IFUPATH90.swl.thr1_state;
thread_status[362] = `IFUPATH90.swl.thr2_state;
thread_status[363] = `IFUPATH90.swl.thr3_state;
thread_status[364] = `IFUPATH91.swl.thr0_state;
thread_status[365] = `IFUPATH91.swl.thr1_state;
thread_status[366] = `IFUPATH91.swl.thr2_state;
thread_status[367] = `IFUPATH91.swl.thr3_state;
thread_status[368] = `IFUPATH92.swl.thr0_state;
thread_status[369] = `IFUPATH92.swl.thr1_state;
thread_status[370] = `IFUPATH92.swl.thr2_state;
thread_status[371] = `IFUPATH92.swl.thr3_state;
thread_status[372] = `IFUPATH93.swl.thr0_state;
thread_status[373] = `IFUPATH93.swl.thr1_state;
thread_status[374] = `IFUPATH93.swl.thr2_state;
thread_status[375] = `IFUPATH93.swl.thr3_state;
thread_status[376] = `IFUPATH94.swl.thr0_state;
thread_status[377] = `IFUPATH94.swl.thr1_state;
thread_status[378] = `IFUPATH94.swl.thr2_state;
thread_status[379] = `IFUPATH94.swl.thr3_state;
thread_status[380] = `IFUPATH95.swl.thr0_state;
thread_status[381] = `IFUPATH95.swl.thr1_state;
thread_status[382] = `IFUPATH95.swl.thr2_state;
thread_status[383] = `IFUPATH95.swl.thr3_state;
thread_status[384] = `IFUPATH96.swl.thr0_state;
thread_status[385] = `IFUPATH96.swl.thr1_state;
thread_status[386] = `IFUPATH96.swl.thr2_state;
thread_status[387] = `IFUPATH96.swl.thr3_state;
thread_status[388] = `IFUPATH97.swl.thr0_state;
thread_status[389] = `IFUPATH97.swl.thr1_state;
thread_status[390] = `IFUPATH97.swl.thr2_state;
thread_status[391] = `IFUPATH97.swl.thr3_state;
thread_status[392] = `IFUPATH98.swl.thr0_state;
thread_status[393] = `IFUPATH98.swl.thr1_state;
thread_status[394] = `IFUPATH98.swl.thr2_state;
thread_status[395] = `IFUPATH98.swl.thr3_state;
thread_status[396] = `IFUPATH99.swl.thr0_state;
thread_status[397] = `IFUPATH99.swl.thr1_state;
thread_status[398] = `IFUPATH99.swl.thr2_state;
thread_status[399] = `IFUPATH99.swl.thr3_state;
thread_status[400] = `IFUPATH100.swl.thr0_state;
thread_status[401] = `IFUPATH100.swl.thr1_state;
thread_status[402] = `IFUPATH100.swl.thr2_state;
thread_status[403] = `IFUPATH100.swl.thr3_state;
thread_status[404] = `IFUPATH101.swl.thr0_state;
thread_status[405] = `IFUPATH101.swl.thr1_state;
thread_status[406] = `IFUPATH101.swl.thr2_state;
thread_status[407] = `IFUPATH101.swl.thr3_state;
thread_status[408] = `IFUPATH102.swl.thr0_state;
thread_status[409] = `IFUPATH102.swl.thr1_state;
thread_status[410] = `IFUPATH102.swl.thr2_state;
thread_status[411] = `IFUPATH102.swl.thr3_state;
thread_status[412] = `IFUPATH103.swl.thr0_state;
thread_status[413] = `IFUPATH103.swl.thr1_state;
thread_status[414] = `IFUPATH103.swl.thr2_state;
thread_status[415] = `IFUPATH103.swl.thr3_state;
thread_status[416] = `IFUPATH104.swl.thr0_state;
thread_status[417] = `IFUPATH104.swl.thr1_state;
thread_status[418] = `IFUPATH104.swl.thr2_state;
thread_status[419] = `IFUPATH104.swl.thr3_state;
thread_status[420] = `IFUPATH105.swl.thr0_state;
thread_status[421] = `IFUPATH105.swl.thr1_state;
thread_status[422] = `IFUPATH105.swl.thr2_state;
thread_status[423] = `IFUPATH105.swl.thr3_state;
thread_status[424] = `IFUPATH106.swl.thr0_state;
thread_status[425] = `IFUPATH106.swl.thr1_state;
thread_status[426] = `IFUPATH106.swl.thr2_state;
thread_status[427] = `IFUPATH106.swl.thr3_state;
thread_status[428] = `IFUPATH107.swl.thr0_state;
thread_status[429] = `IFUPATH107.swl.thr1_state;
thread_status[430] = `IFUPATH107.swl.thr2_state;
thread_status[431] = `IFUPATH107.swl.thr3_state;
thread_status[432] = `IFUPATH108.swl.thr0_state;
thread_status[433] = `IFUPATH108.swl.thr1_state;
thread_status[434] = `IFUPATH108.swl.thr2_state;
thread_status[435] = `IFUPATH108.swl.thr3_state;
thread_status[436] = `IFUPATH109.swl.thr0_state;
thread_status[437] = `IFUPATH109.swl.thr1_state;
thread_status[438] = `IFUPATH109.swl.thr2_state;
thread_status[439] = `IFUPATH109.swl.thr3_state;
thread_status[440] = `IFUPATH110.swl.thr0_state;
thread_status[441] = `IFUPATH110.swl.thr1_state;
thread_status[442] = `IFUPATH110.swl.thr2_state;
thread_status[443] = `IFUPATH110.swl.thr3_state;
thread_status[444] = `IFUPATH111.swl.thr0_state;
thread_status[445] = `IFUPATH111.swl.thr1_state;
thread_status[446] = `IFUPATH111.swl.thr2_state;
thread_status[447] = `IFUPATH111.swl.thr3_state;
thread_status[448] = `IFUPATH112.swl.thr0_state;
thread_status[449] = `IFUPATH112.swl.thr1_state;
thread_status[450] = `IFUPATH112.swl.thr2_state;
thread_status[451] = `IFUPATH112.swl.thr3_state;
thread_status[452] = `IFUPATH113.swl.thr0_state;
thread_status[453] = `IFUPATH113.swl.thr1_state;
thread_status[454] = `IFUPATH113.swl.thr2_state;
thread_status[455] = `IFUPATH113.swl.thr3_state;
thread_status[456] = `IFUPATH114.swl.thr0_state;
thread_status[457] = `IFUPATH114.swl.thr1_state;
thread_status[458] = `IFUPATH114.swl.thr2_state;
thread_status[459] = `IFUPATH114.swl.thr3_state;
thread_status[460] = `IFUPATH115.swl.thr0_state;
thread_status[461] = `IFUPATH115.swl.thr1_state;
thread_status[462] = `IFUPATH115.swl.thr2_state;
thread_status[463] = `IFUPATH115.swl.thr3_state;
thread_status[464] = `IFUPATH116.swl.thr0_state;
thread_status[465] = `IFUPATH116.swl.thr1_state;
thread_status[466] = `IFUPATH116.swl.thr2_state;
thread_status[467] = `IFUPATH116.swl.thr3_state;
thread_status[468] = `IFUPATH117.swl.thr0_state;
thread_status[469] = `IFUPATH117.swl.thr1_state;
thread_status[470] = `IFUPATH117.swl.thr2_state;
thread_status[471] = `IFUPATH117.swl.thr3_state;
thread_status[472] = `IFUPATH118.swl.thr0_state;
thread_status[473] = `IFUPATH118.swl.thr1_state;
thread_status[474] = `IFUPATH118.swl.thr2_state;
thread_status[475] = `IFUPATH118.swl.thr3_state;
thread_status[476] = `IFUPATH119.swl.thr0_state;
thread_status[477] = `IFUPATH119.swl.thr1_state;
thread_status[478] = `IFUPATH119.swl.thr2_state;
thread_status[479] = `IFUPATH119.swl.thr3_state;
thread_status[480] = `IFUPATH120.swl.thr0_state;
thread_status[481] = `IFUPATH120.swl.thr1_state;
thread_status[482] = `IFUPATH120.swl.thr2_state;
thread_status[483] = `IFUPATH120.swl.thr3_state;
thread_status[484] = `IFUPATH121.swl.thr0_state;
thread_status[485] = `IFUPATH121.swl.thr1_state;
thread_status[486] = `IFUPATH121.swl.thr2_state;
thread_status[487] = `IFUPATH121.swl.thr3_state;
thread_status[488] = `IFUPATH122.swl.thr0_state;
thread_status[489] = `IFUPATH122.swl.thr1_state;
thread_status[490] = `IFUPATH122.swl.thr2_state;
thread_status[491] = `IFUPATH122.swl.thr3_state;
thread_status[492] = `IFUPATH123.swl.thr0_state;
thread_status[493] = `IFUPATH123.swl.thr1_state;
thread_status[494] = `IFUPATH123.swl.thr2_state;
thread_status[495] = `IFUPATH123.swl.thr3_state;
thread_status[496] = `IFUPATH124.swl.thr0_state;
thread_status[497] = `IFUPATH124.swl.thr1_state;
thread_status[498] = `IFUPATH124.swl.thr2_state;
thread_status[499] = `IFUPATH124.swl.thr3_state;
thread_status[500] = `IFUPATH125.swl.thr0_state;
thread_status[501] = `IFUPATH125.swl.thr1_state;
thread_status[502] = `IFUPATH125.swl.thr2_state;
thread_status[503] = `IFUPATH125.swl.thr3_state;
thread_status[504] = `IFUPATH126.swl.thr0_state;
thread_status[505] = `IFUPATH126.swl.thr1_state;
thread_status[506] = `IFUPATH126.swl.thr2_state;
thread_status[507] = `IFUPATH126.swl.thr3_state;
thread_status[508] = `IFUPATH127.swl.thr0_state;
thread_status[509] = `IFUPATH127.swl.thr1_state;
thread_status[510] = `IFUPATH127.swl.thr2_state;
thread_status[511] = `IFUPATH127.swl.thr3_state;
thread_status[512] = `IFUPATH128.swl.thr0_state;
thread_status[513] = `IFUPATH128.swl.thr1_state;
thread_status[514] = `IFUPATH128.swl.thr2_state;
thread_status[515] = `IFUPATH128.swl.thr3_state;
thread_status[516] = `IFUPATH129.swl.thr0_state;
thread_status[517] = `IFUPATH129.swl.thr1_state;
thread_status[518] = `IFUPATH129.swl.thr2_state;
thread_status[519] = `IFUPATH129.swl.thr3_state;
thread_status[520] = `IFUPATH130.swl.thr0_state;
thread_status[521] = `IFUPATH130.swl.thr1_state;
thread_status[522] = `IFUPATH130.swl.thr2_state;
thread_status[523] = `IFUPATH130.swl.thr3_state;
thread_status[524] = `IFUPATH131.swl.thr0_state;
thread_status[525] = `IFUPATH131.swl.thr1_state;
thread_status[526] = `IFUPATH131.swl.thr2_state;
thread_status[527] = `IFUPATH131.swl.thr3_state;
thread_status[528] = `IFUPATH132.swl.thr0_state;
thread_status[529] = `IFUPATH132.swl.thr1_state;
thread_status[530] = `IFUPATH132.swl.thr2_state;
thread_status[531] = `IFUPATH132.swl.thr3_state;
thread_status[532] = `IFUPATH133.swl.thr0_state;
thread_status[533] = `IFUPATH133.swl.thr1_state;
thread_status[534] = `IFUPATH133.swl.thr2_state;
thread_status[535] = `IFUPATH133.swl.thr3_state;
thread_status[536] = `IFUPATH134.swl.thr0_state;
thread_status[537] = `IFUPATH134.swl.thr1_state;
thread_status[538] = `IFUPATH134.swl.thr2_state;
thread_status[539] = `IFUPATH134.swl.thr3_state;
thread_status[540] = `IFUPATH135.swl.thr0_state;
thread_status[541] = `IFUPATH135.swl.thr1_state;
thread_status[542] = `IFUPATH135.swl.thr2_state;
thread_status[543] = `IFUPATH135.swl.thr3_state;
thread_status[544] = `IFUPATH136.swl.thr0_state;
thread_status[545] = `IFUPATH136.swl.thr1_state;
thread_status[546] = `IFUPATH136.swl.thr2_state;
thread_status[547] = `IFUPATH136.swl.thr3_state;
thread_status[548] = `IFUPATH137.swl.thr0_state;
thread_status[549] = `IFUPATH137.swl.thr1_state;
thread_status[550] = `IFUPATH137.swl.thr2_state;
thread_status[551] = `IFUPATH137.swl.thr3_state;
thread_status[552] = `IFUPATH138.swl.thr0_state;
thread_status[553] = `IFUPATH138.swl.thr1_state;
thread_status[554] = `IFUPATH138.swl.thr2_state;
thread_status[555] = `IFUPATH138.swl.thr3_state;
thread_status[556] = `IFUPATH139.swl.thr0_state;
thread_status[557] = `IFUPATH139.swl.thr1_state;
thread_status[558] = `IFUPATH139.swl.thr2_state;
thread_status[559] = `IFUPATH139.swl.thr3_state;
thread_status[560] = `IFUPATH140.swl.thr0_state;
thread_status[561] = `IFUPATH140.swl.thr1_state;
thread_status[562] = `IFUPATH140.swl.thr2_state;
thread_status[563] = `IFUPATH140.swl.thr3_state;
thread_status[564] = `IFUPATH141.swl.thr0_state;
thread_status[565] = `IFUPATH141.swl.thr1_state;
thread_status[566] = `IFUPATH141.swl.thr2_state;
thread_status[567] = `IFUPATH141.swl.thr3_state;
thread_status[568] = `IFUPATH142.swl.thr0_state;
thread_status[569] = `IFUPATH142.swl.thr1_state;
thread_status[570] = `IFUPATH142.swl.thr2_state;
thread_status[571] = `IFUPATH142.swl.thr3_state;
thread_status[572] = `IFUPATH143.swl.thr0_state;
thread_status[573] = `IFUPATH143.swl.thr1_state;
thread_status[574] = `IFUPATH143.swl.thr2_state;
thread_status[575] = `IFUPATH143.swl.thr3_state;
thread_status[576] = `IFUPATH144.swl.thr0_state;
thread_status[577] = `IFUPATH144.swl.thr1_state;
thread_status[578] = `IFUPATH144.swl.thr2_state;
thread_status[579] = `IFUPATH144.swl.thr3_state;
thread_status[580] = `IFUPATH145.swl.thr0_state;
thread_status[581] = `IFUPATH145.swl.thr1_state;
thread_status[582] = `IFUPATH145.swl.thr2_state;
thread_status[583] = `IFUPATH145.swl.thr3_state;
thread_status[584] = `IFUPATH146.swl.thr0_state;
thread_status[585] = `IFUPATH146.swl.thr1_state;
thread_status[586] = `IFUPATH146.swl.thr2_state;
thread_status[587] = `IFUPATH146.swl.thr3_state;
thread_status[588] = `IFUPATH147.swl.thr0_state;
thread_status[589] = `IFUPATH147.swl.thr1_state;
thread_status[590] = `IFUPATH147.swl.thr2_state;
thread_status[591] = `IFUPATH147.swl.thr3_state;
thread_status[592] = `IFUPATH148.swl.thr0_state;
thread_status[593] = `IFUPATH148.swl.thr1_state;
thread_status[594] = `IFUPATH148.swl.thr2_state;
thread_status[595] = `IFUPATH148.swl.thr3_state;
thread_status[596] = `IFUPATH149.swl.thr0_state;
thread_status[597] = `IFUPATH149.swl.thr1_state;
thread_status[598] = `IFUPATH149.swl.thr2_state;
thread_status[599] = `IFUPATH149.swl.thr3_state;
thread_status[600] = `IFUPATH150.swl.thr0_state;
thread_status[601] = `IFUPATH150.swl.thr1_state;
thread_status[602] = `IFUPATH150.swl.thr2_state;
thread_status[603] = `IFUPATH150.swl.thr3_state;
thread_status[604] = `IFUPATH151.swl.thr0_state;
thread_status[605] = `IFUPATH151.swl.thr1_state;
thread_status[606] = `IFUPATH151.swl.thr2_state;
thread_status[607] = `IFUPATH151.swl.thr3_state;
thread_status[608] = `IFUPATH152.swl.thr0_state;
thread_status[609] = `IFUPATH152.swl.thr1_state;
thread_status[610] = `IFUPATH152.swl.thr2_state;
thread_status[611] = `IFUPATH152.swl.thr3_state;
thread_status[612] = `IFUPATH153.swl.thr0_state;
thread_status[613] = `IFUPATH153.swl.thr1_state;
thread_status[614] = `IFUPATH153.swl.thr2_state;
thread_status[615] = `IFUPATH153.swl.thr3_state;
thread_status[616] = `IFUPATH154.swl.thr0_state;
thread_status[617] = `IFUPATH154.swl.thr1_state;
thread_status[618] = `IFUPATH154.swl.thr2_state;
thread_status[619] = `IFUPATH154.swl.thr3_state;
thread_status[620] = `IFUPATH155.swl.thr0_state;
thread_status[621] = `IFUPATH155.swl.thr1_state;
thread_status[622] = `IFUPATH155.swl.thr2_state;
thread_status[623] = `IFUPATH155.swl.thr3_state;
thread_status[624] = `IFUPATH156.swl.thr0_state;
thread_status[625] = `IFUPATH156.swl.thr1_state;
thread_status[626] = `IFUPATH156.swl.thr2_state;
thread_status[627] = `IFUPATH156.swl.thr3_state;
thread_status[628] = `IFUPATH157.swl.thr0_state;
thread_status[629] = `IFUPATH157.swl.thr1_state;
thread_status[630] = `IFUPATH157.swl.thr2_state;
thread_status[631] = `IFUPATH157.swl.thr3_state;
thread_status[632] = `IFUPATH158.swl.thr0_state;
thread_status[633] = `IFUPATH158.swl.thr1_state;
thread_status[634] = `IFUPATH158.swl.thr2_state;
thread_status[635] = `IFUPATH158.swl.thr3_state;
thread_status[636] = `IFUPATH159.swl.thr0_state;
thread_status[637] = `IFUPATH159.swl.thr1_state;
thread_status[638] = `IFUPATH159.swl.thr2_state;
thread_status[639] = `IFUPATH159.swl.thr3_state;
thread_status[640] = `IFUPATH160.swl.thr0_state;
thread_status[641] = `IFUPATH160.swl.thr1_state;
thread_status[642] = `IFUPATH160.swl.thr2_state;
thread_status[643] = `IFUPATH160.swl.thr3_state;
thread_status[644] = `IFUPATH161.swl.thr0_state;
thread_status[645] = `IFUPATH161.swl.thr1_state;
thread_status[646] = `IFUPATH161.swl.thr2_state;
thread_status[647] = `IFUPATH161.swl.thr3_state;
thread_status[648] = `IFUPATH162.swl.thr0_state;
thread_status[649] = `IFUPATH162.swl.thr1_state;
thread_status[650] = `IFUPATH162.swl.thr2_state;
thread_status[651] = `IFUPATH162.swl.thr3_state;
thread_status[652] = `IFUPATH163.swl.thr0_state;
thread_status[653] = `IFUPATH163.swl.thr1_state;
thread_status[654] = `IFUPATH163.swl.thr2_state;
thread_status[655] = `IFUPATH163.swl.thr3_state;
thread_status[656] = `IFUPATH164.swl.thr0_state;
thread_status[657] = `IFUPATH164.swl.thr1_state;
thread_status[658] = `IFUPATH164.swl.thr2_state;
thread_status[659] = `IFUPATH164.swl.thr3_state;
thread_status[660] = `IFUPATH165.swl.thr0_state;
thread_status[661] = `IFUPATH165.swl.thr1_state;
thread_status[662] = `IFUPATH165.swl.thr2_state;
thread_status[663] = `IFUPATH165.swl.thr3_state;
thread_status[664] = `IFUPATH166.swl.thr0_state;
thread_status[665] = `IFUPATH166.swl.thr1_state;
thread_status[666] = `IFUPATH166.swl.thr2_state;
thread_status[667] = `IFUPATH166.swl.thr3_state;
thread_status[668] = `IFUPATH167.swl.thr0_state;
thread_status[669] = `IFUPATH167.swl.thr1_state;
thread_status[670] = `IFUPATH167.swl.thr2_state;
thread_status[671] = `IFUPATH167.swl.thr3_state;
thread_status[672] = `IFUPATH168.swl.thr0_state;
thread_status[673] = `IFUPATH168.swl.thr1_state;
thread_status[674] = `IFUPATH168.swl.thr2_state;
thread_status[675] = `IFUPATH168.swl.thr3_state;
thread_status[676] = `IFUPATH169.swl.thr0_state;
thread_status[677] = `IFUPATH169.swl.thr1_state;
thread_status[678] = `IFUPATH169.swl.thr2_state;
thread_status[679] = `IFUPATH169.swl.thr3_state;
thread_status[680] = `IFUPATH170.swl.thr0_state;
thread_status[681] = `IFUPATH170.swl.thr1_state;
thread_status[682] = `IFUPATH170.swl.thr2_state;
thread_status[683] = `IFUPATH170.swl.thr3_state;
thread_status[684] = `IFUPATH171.swl.thr0_state;
thread_status[685] = `IFUPATH171.swl.thr1_state;
thread_status[686] = `IFUPATH171.swl.thr2_state;
thread_status[687] = `IFUPATH171.swl.thr3_state;
thread_status[688] = `IFUPATH172.swl.thr0_state;
thread_status[689] = `IFUPATH172.swl.thr1_state;
thread_status[690] = `IFUPATH172.swl.thr2_state;
thread_status[691] = `IFUPATH172.swl.thr3_state;
thread_status[692] = `IFUPATH173.swl.thr0_state;
thread_status[693] = `IFUPATH173.swl.thr1_state;
thread_status[694] = `IFUPATH173.swl.thr2_state;
thread_status[695] = `IFUPATH173.swl.thr3_state;
thread_status[696] = `IFUPATH174.swl.thr0_state;
thread_status[697] = `IFUPATH174.swl.thr1_state;
thread_status[698] = `IFUPATH174.swl.thr2_state;
thread_status[699] = `IFUPATH174.swl.thr3_state;
thread_status[700] = `IFUPATH175.swl.thr0_state;
thread_status[701] = `IFUPATH175.swl.thr1_state;
thread_status[702] = `IFUPATH175.swl.thr2_state;
thread_status[703] = `IFUPATH175.swl.thr3_state;
thread_status[704] = `IFUPATH176.swl.thr0_state;
thread_status[705] = `IFUPATH176.swl.thr1_state;
thread_status[706] = `IFUPATH176.swl.thr2_state;
thread_status[707] = `IFUPATH176.swl.thr3_state;
thread_status[708] = `IFUPATH177.swl.thr0_state;
thread_status[709] = `IFUPATH177.swl.thr1_state;
thread_status[710] = `IFUPATH177.swl.thr2_state;
thread_status[711] = `IFUPATH177.swl.thr3_state;
thread_status[712] = `IFUPATH178.swl.thr0_state;
thread_status[713] = `IFUPATH178.swl.thr1_state;
thread_status[714] = `IFUPATH178.swl.thr2_state;
thread_status[715] = `IFUPATH178.swl.thr3_state;
thread_status[716] = `IFUPATH179.swl.thr0_state;
thread_status[717] = `IFUPATH179.swl.thr1_state;
thread_status[718] = `IFUPATH179.swl.thr2_state;
thread_status[719] = `IFUPATH179.swl.thr3_state;
thread_status[720] = `IFUPATH180.swl.thr0_state;
thread_status[721] = `IFUPATH180.swl.thr1_state;
thread_status[722] = `IFUPATH180.swl.thr2_state;
thread_status[723] = `IFUPATH180.swl.thr3_state;
thread_status[724] = `IFUPATH181.swl.thr0_state;
thread_status[725] = `IFUPATH181.swl.thr1_state;
thread_status[726] = `IFUPATH181.swl.thr2_state;
thread_status[727] = `IFUPATH181.swl.thr3_state;
thread_status[728] = `IFUPATH182.swl.thr0_state;
thread_status[729] = `IFUPATH182.swl.thr1_state;
thread_status[730] = `IFUPATH182.swl.thr2_state;
thread_status[731] = `IFUPATH182.swl.thr3_state;
thread_status[732] = `IFUPATH183.swl.thr0_state;
thread_status[733] = `IFUPATH183.swl.thr1_state;
thread_status[734] = `IFUPATH183.swl.thr2_state;
thread_status[735] = `IFUPATH183.swl.thr3_state;
thread_status[736] = `IFUPATH184.swl.thr0_state;
thread_status[737] = `IFUPATH184.swl.thr1_state;
thread_status[738] = `IFUPATH184.swl.thr2_state;
thread_status[739] = `IFUPATH184.swl.thr3_state;
thread_status[740] = `IFUPATH185.swl.thr0_state;
thread_status[741] = `IFUPATH185.swl.thr1_state;
thread_status[742] = `IFUPATH185.swl.thr2_state;
thread_status[743] = `IFUPATH185.swl.thr3_state;
thread_status[744] = `IFUPATH186.swl.thr0_state;
thread_status[745] = `IFUPATH186.swl.thr1_state;
thread_status[746] = `IFUPATH186.swl.thr2_state;
thread_status[747] = `IFUPATH186.swl.thr3_state;
thread_status[748] = `IFUPATH187.swl.thr0_state;
thread_status[749] = `IFUPATH187.swl.thr1_state;
thread_status[750] = `IFUPATH187.swl.thr2_state;
thread_status[751] = `IFUPATH187.swl.thr3_state;
thread_status[752] = `IFUPATH188.swl.thr0_state;
thread_status[753] = `IFUPATH188.swl.thr1_state;
thread_status[754] = `IFUPATH188.swl.thr2_state;
thread_status[755] = `IFUPATH188.swl.thr3_state;
thread_status[756] = `IFUPATH189.swl.thr0_state;
thread_status[757] = `IFUPATH189.swl.thr1_state;
thread_status[758] = `IFUPATH189.swl.thr2_state;
thread_status[759] = `IFUPATH189.swl.thr3_state;
thread_status[760] = `IFUPATH190.swl.thr0_state;
thread_status[761] = `IFUPATH190.swl.thr1_state;
thread_status[762] = `IFUPATH190.swl.thr2_state;
thread_status[763] = `IFUPATH190.swl.thr3_state;
thread_status[764] = `IFUPATH191.swl.thr0_state;
thread_status[765] = `IFUPATH191.swl.thr1_state;
thread_status[766] = `IFUPATH191.swl.thr2_state;
thread_status[767] = `IFUPATH191.swl.thr3_state;
thread_status[768] = `IFUPATH192.swl.thr0_state;
thread_status[769] = `IFUPATH192.swl.thr1_state;
thread_status[770] = `IFUPATH192.swl.thr2_state;
thread_status[771] = `IFUPATH192.swl.thr3_state;
thread_status[772] = `IFUPATH193.swl.thr0_state;
thread_status[773] = `IFUPATH193.swl.thr1_state;
thread_status[774] = `IFUPATH193.swl.thr2_state;
thread_status[775] = `IFUPATH193.swl.thr3_state;
thread_status[776] = `IFUPATH194.swl.thr0_state;
thread_status[777] = `IFUPATH194.swl.thr1_state;
thread_status[778] = `IFUPATH194.swl.thr2_state;
thread_status[779] = `IFUPATH194.swl.thr3_state;
thread_status[780] = `IFUPATH195.swl.thr0_state;
thread_status[781] = `IFUPATH195.swl.thr1_state;
thread_status[782] = `IFUPATH195.swl.thr2_state;
thread_status[783] = `IFUPATH195.swl.thr3_state;
thread_status[784] = `IFUPATH196.swl.thr0_state;
thread_status[785] = `IFUPATH196.swl.thr1_state;
thread_status[786] = `IFUPATH196.swl.thr2_state;
thread_status[787] = `IFUPATH196.swl.thr3_state;
thread_status[788] = `IFUPATH197.swl.thr0_state;
thread_status[789] = `IFUPATH197.swl.thr1_state;
thread_status[790] = `IFUPATH197.swl.thr2_state;
thread_status[791] = `IFUPATH197.swl.thr3_state;
thread_status[792] = `IFUPATH198.swl.thr0_state;
thread_status[793] = `IFUPATH198.swl.thr1_state;
thread_status[794] = `IFUPATH198.swl.thr2_state;
thread_status[795] = `IFUPATH198.swl.thr3_state;
thread_status[796] = `IFUPATH199.swl.thr0_state;
thread_status[797] = `IFUPATH199.swl.thr1_state;
thread_status[798] = `IFUPATH199.swl.thr2_state;
thread_status[799] = `IFUPATH199.swl.thr3_state;
thread_status[800] = `IFUPATH200.swl.thr0_state;
thread_status[801] = `IFUPATH200.swl.thr1_state;
thread_status[802] = `IFUPATH200.swl.thr2_state;
thread_status[803] = `IFUPATH200.swl.thr3_state;
thread_status[804] = `IFUPATH201.swl.thr0_state;
thread_status[805] = `IFUPATH201.swl.thr1_state;
thread_status[806] = `IFUPATH201.swl.thr2_state;
thread_status[807] = `IFUPATH201.swl.thr3_state;
thread_status[808] = `IFUPATH202.swl.thr0_state;
thread_status[809] = `IFUPATH202.swl.thr1_state;
thread_status[810] = `IFUPATH202.swl.thr2_state;
thread_status[811] = `IFUPATH202.swl.thr3_state;
thread_status[812] = `IFUPATH203.swl.thr0_state;
thread_status[813] = `IFUPATH203.swl.thr1_state;
thread_status[814] = `IFUPATH203.swl.thr2_state;
thread_status[815] = `IFUPATH203.swl.thr3_state;
thread_status[816] = `IFUPATH204.swl.thr0_state;
thread_status[817] = `IFUPATH204.swl.thr1_state;
thread_status[818] = `IFUPATH204.swl.thr2_state;
thread_status[819] = `IFUPATH204.swl.thr3_state;
thread_status[820] = `IFUPATH205.swl.thr0_state;
thread_status[821] = `IFUPATH205.swl.thr1_state;
thread_status[822] = `IFUPATH205.swl.thr2_state;
thread_status[823] = `IFUPATH205.swl.thr3_state;
thread_status[824] = `IFUPATH206.swl.thr0_state;
thread_status[825] = `IFUPATH206.swl.thr1_state;
thread_status[826] = `IFUPATH206.swl.thr2_state;
thread_status[827] = `IFUPATH206.swl.thr3_state;
thread_status[828] = `IFUPATH207.swl.thr0_state;
thread_status[829] = `IFUPATH207.swl.thr1_state;
thread_status[830] = `IFUPATH207.swl.thr2_state;
thread_status[831] = `IFUPATH207.swl.thr3_state;
thread_status[832] = `IFUPATH208.swl.thr0_state;
thread_status[833] = `IFUPATH208.swl.thr1_state;
thread_status[834] = `IFUPATH208.swl.thr2_state;
thread_status[835] = `IFUPATH208.swl.thr3_state;
thread_status[836] = `IFUPATH209.swl.thr0_state;
thread_status[837] = `IFUPATH209.swl.thr1_state;
thread_status[838] = `IFUPATH209.swl.thr2_state;
thread_status[839] = `IFUPATH209.swl.thr3_state;
thread_status[840] = `IFUPATH210.swl.thr0_state;
thread_status[841] = `IFUPATH210.swl.thr1_state;
thread_status[842] = `IFUPATH210.swl.thr2_state;
thread_status[843] = `IFUPATH210.swl.thr3_state;
thread_status[844] = `IFUPATH211.swl.thr0_state;
thread_status[845] = `IFUPATH211.swl.thr1_state;
thread_status[846] = `IFUPATH211.swl.thr2_state;
thread_status[847] = `IFUPATH211.swl.thr3_state;
thread_status[848] = `IFUPATH212.swl.thr0_state;
thread_status[849] = `IFUPATH212.swl.thr1_state;
thread_status[850] = `IFUPATH212.swl.thr2_state;
thread_status[851] = `IFUPATH212.swl.thr3_state;
thread_status[852] = `IFUPATH213.swl.thr0_state;
thread_status[853] = `IFUPATH213.swl.thr1_state;
thread_status[854] = `IFUPATH213.swl.thr2_state;
thread_status[855] = `IFUPATH213.swl.thr3_state;
thread_status[856] = `IFUPATH214.swl.thr0_state;
thread_status[857] = `IFUPATH214.swl.thr1_state;
thread_status[858] = `IFUPATH214.swl.thr2_state;
thread_status[859] = `IFUPATH214.swl.thr3_state;
thread_status[860] = `IFUPATH215.swl.thr0_state;
thread_status[861] = `IFUPATH215.swl.thr1_state;
thread_status[862] = `IFUPATH215.swl.thr2_state;
thread_status[863] = `IFUPATH215.swl.thr3_state;
thread_status[864] = `IFUPATH216.swl.thr0_state;
thread_status[865] = `IFUPATH216.swl.thr1_state;
thread_status[866] = `IFUPATH216.swl.thr2_state;
thread_status[867] = `IFUPATH216.swl.thr3_state;
thread_status[868] = `IFUPATH217.swl.thr0_state;
thread_status[869] = `IFUPATH217.swl.thr1_state;
thread_status[870] = `IFUPATH217.swl.thr2_state;
thread_status[871] = `IFUPATH217.swl.thr3_state;
thread_status[872] = `IFUPATH218.swl.thr0_state;
thread_status[873] = `IFUPATH218.swl.thr1_state;
thread_status[874] = `IFUPATH218.swl.thr2_state;
thread_status[875] = `IFUPATH218.swl.thr3_state;
thread_status[876] = `IFUPATH219.swl.thr0_state;
thread_status[877] = `IFUPATH219.swl.thr1_state;
thread_status[878] = `IFUPATH219.swl.thr2_state;
thread_status[879] = `IFUPATH219.swl.thr3_state;
thread_status[880] = `IFUPATH220.swl.thr0_state;
thread_status[881] = `IFUPATH220.swl.thr1_state;
thread_status[882] = `IFUPATH220.swl.thr2_state;
thread_status[883] = `IFUPATH220.swl.thr3_state;
thread_status[884] = `IFUPATH221.swl.thr0_state;
thread_status[885] = `IFUPATH221.swl.thr1_state;
thread_status[886] = `IFUPATH221.swl.thr2_state;
thread_status[887] = `IFUPATH221.swl.thr3_state;
thread_status[888] = `IFUPATH222.swl.thr0_state;
thread_status[889] = `IFUPATH222.swl.thr1_state;
thread_status[890] = `IFUPATH222.swl.thr2_state;
thread_status[891] = `IFUPATH222.swl.thr3_state;
thread_status[892] = `IFUPATH223.swl.thr0_state;
thread_status[893] = `IFUPATH223.swl.thr1_state;
thread_status[894] = `IFUPATH223.swl.thr2_state;
thread_status[895] = `IFUPATH223.swl.thr3_state;
thread_status[896] = `IFUPATH224.swl.thr0_state;
thread_status[897] = `IFUPATH224.swl.thr1_state;
thread_status[898] = `IFUPATH224.swl.thr2_state;
thread_status[899] = `IFUPATH224.swl.thr3_state;
thread_status[900] = `IFUPATH225.swl.thr0_state;
thread_status[901] = `IFUPATH225.swl.thr1_state;
thread_status[902] = `IFUPATH225.swl.thr2_state;
thread_status[903] = `IFUPATH225.swl.thr3_state;
thread_status[904] = `IFUPATH226.swl.thr0_state;
thread_status[905] = `IFUPATH226.swl.thr1_state;
thread_status[906] = `IFUPATH226.swl.thr2_state;
thread_status[907] = `IFUPATH226.swl.thr3_state;
thread_status[908] = `IFUPATH227.swl.thr0_state;
thread_status[909] = `IFUPATH227.swl.thr1_state;
thread_status[910] = `IFUPATH227.swl.thr2_state;
thread_status[911] = `IFUPATH227.swl.thr3_state;
thread_status[912] = `IFUPATH228.swl.thr0_state;
thread_status[913] = `IFUPATH228.swl.thr1_state;
thread_status[914] = `IFUPATH228.swl.thr2_state;
thread_status[915] = `IFUPATH228.swl.thr3_state;
thread_status[916] = `IFUPATH229.swl.thr0_state;
thread_status[917] = `IFUPATH229.swl.thr1_state;
thread_status[918] = `IFUPATH229.swl.thr2_state;
thread_status[919] = `IFUPATH229.swl.thr3_state;
thread_status[920] = `IFUPATH230.swl.thr0_state;
thread_status[921] = `IFUPATH230.swl.thr1_state;
thread_status[922] = `IFUPATH230.swl.thr2_state;
thread_status[923] = `IFUPATH230.swl.thr3_state;
thread_status[924] = `IFUPATH231.swl.thr0_state;
thread_status[925] = `IFUPATH231.swl.thr1_state;
thread_status[926] = `IFUPATH231.swl.thr2_state;
thread_status[927] = `IFUPATH231.swl.thr3_state;
thread_status[928] = `IFUPATH232.swl.thr0_state;
thread_status[929] = `IFUPATH232.swl.thr1_state;
thread_status[930] = `IFUPATH232.swl.thr2_state;
thread_status[931] = `IFUPATH232.swl.thr3_state;
thread_status[932] = `IFUPATH233.swl.thr0_state;
thread_status[933] = `IFUPATH233.swl.thr1_state;
thread_status[934] = `IFUPATH233.swl.thr2_state;
thread_status[935] = `IFUPATH233.swl.thr3_state;
thread_status[936] = `IFUPATH234.swl.thr0_state;
thread_status[937] = `IFUPATH234.swl.thr1_state;
thread_status[938] = `IFUPATH234.swl.thr2_state;
thread_status[939] = `IFUPATH234.swl.thr3_state;
thread_status[940] = `IFUPATH235.swl.thr0_state;
thread_status[941] = `IFUPATH235.swl.thr1_state;
thread_status[942] = `IFUPATH235.swl.thr2_state;
thread_status[943] = `IFUPATH235.swl.thr3_state;
thread_status[944] = `IFUPATH236.swl.thr0_state;
thread_status[945] = `IFUPATH236.swl.thr1_state;
thread_status[946] = `IFUPATH236.swl.thr2_state;
thread_status[947] = `IFUPATH236.swl.thr3_state;
thread_status[948] = `IFUPATH237.swl.thr0_state;
thread_status[949] = `IFUPATH237.swl.thr1_state;
thread_status[950] = `IFUPATH237.swl.thr2_state;
thread_status[951] = `IFUPATH237.swl.thr3_state;
thread_status[952] = `IFUPATH238.swl.thr0_state;
thread_status[953] = `IFUPATH238.swl.thr1_state;
thread_status[954] = `IFUPATH238.swl.thr2_state;
thread_status[955] = `IFUPATH238.swl.thr3_state;
thread_status[956] = `IFUPATH239.swl.thr0_state;
thread_status[957] = `IFUPATH239.swl.thr1_state;
thread_status[958] = `IFUPATH239.swl.thr2_state;
thread_status[959] = `IFUPATH239.swl.thr3_state;
thread_status[960] = `IFUPATH240.swl.thr0_state;
thread_status[961] = `IFUPATH240.swl.thr1_state;
thread_status[962] = `IFUPATH240.swl.thr2_state;
thread_status[963] = `IFUPATH240.swl.thr3_state;
thread_status[964] = `IFUPATH241.swl.thr0_state;
thread_status[965] = `IFUPATH241.swl.thr1_state;
thread_status[966] = `IFUPATH241.swl.thr2_state;
thread_status[967] = `IFUPATH241.swl.thr3_state;
thread_status[968] = `IFUPATH242.swl.thr0_state;
thread_status[969] = `IFUPATH242.swl.thr1_state;
thread_status[970] = `IFUPATH242.swl.thr2_state;
thread_status[971] = `IFUPATH242.swl.thr3_state;
thread_status[972] = `IFUPATH243.swl.thr0_state;
thread_status[973] = `IFUPATH243.swl.thr1_state;
thread_status[974] = `IFUPATH243.swl.thr2_state;
thread_status[975] = `IFUPATH243.swl.thr3_state;
thread_status[976] = `IFUPATH244.swl.thr0_state;
thread_status[977] = `IFUPATH244.swl.thr1_state;
thread_status[978] = `IFUPATH244.swl.thr2_state;
thread_status[979] = `IFUPATH244.swl.thr3_state;
thread_status[980] = `IFUPATH245.swl.thr0_state;
thread_status[981] = `IFUPATH245.swl.thr1_state;
thread_status[982] = `IFUPATH245.swl.thr2_state;
thread_status[983] = `IFUPATH245.swl.thr3_state;
thread_status[984] = `IFUPATH246.swl.thr0_state;
thread_status[985] = `IFUPATH246.swl.thr1_state;
thread_status[986] = `IFUPATH246.swl.thr2_state;
thread_status[987] = `IFUPATH246.swl.thr3_state;
thread_status[988] = `IFUPATH247.swl.thr0_state;
thread_status[989] = `IFUPATH247.swl.thr1_state;
thread_status[990] = `IFUPATH247.swl.thr2_state;
thread_status[991] = `IFUPATH247.swl.thr3_state;
thread_status[992] = `IFUPATH248.swl.thr0_state;
thread_status[993] = `IFUPATH248.swl.thr1_state;
thread_status[994] = `IFUPATH248.swl.thr2_state;
thread_status[995] = `IFUPATH248.swl.thr3_state;
thread_status[996] = `IFUPATH249.swl.thr0_state;
thread_status[997] = `IFUPATH249.swl.thr1_state;
thread_status[998] = `IFUPATH249.swl.thr2_state;
thread_status[999] = `IFUPATH249.swl.thr3_state;
thread_status[1000] = `IFUPATH250.swl.thr0_state;
thread_status[1001] = `IFUPATH250.swl.thr1_state;
thread_status[1002] = `IFUPATH250.swl.thr2_state;
thread_status[1003] = `IFUPATH250.swl.thr3_state;
thread_status[1004] = `IFUPATH251.swl.thr0_state;
thread_status[1005] = `IFUPATH251.swl.thr1_state;
thread_status[1006] = `IFUPATH251.swl.thr2_state;
thread_status[1007] = `IFUPATH251.swl.thr3_state;
thread_status[1008] = `IFUPATH252.swl.thr0_state;
thread_status[1009] = `IFUPATH252.swl.thr1_state;
thread_status[1010] = `IFUPATH252.swl.thr2_state;
thread_status[1011] = `IFUPATH252.swl.thr3_state;
thread_status[1012] = `IFUPATH253.swl.thr0_state;
thread_status[1013] = `IFUPATH253.swl.thr1_state;
thread_status[1014] = `IFUPATH253.swl.thr2_state;
thread_status[1015] = `IFUPATH253.swl.thr3_state;
thread_status[1016] = `IFUPATH254.swl.thr0_state;
thread_status[1017] = `IFUPATH254.swl.thr1_state;
thread_status[1018] = `IFUPATH254.swl.thr2_state;
thread_status[1019] = `IFUPATH254.swl.thr3_state;
thread_status[1020] = `IFUPATH255.swl.thr0_state;
thread_status[1021] = `IFUPATH255.swl.thr1_state;
thread_status[1022] = `IFUPATH255.swl.thr2_state;
thread_status[1023] = `IFUPATH255.swl.thr3_state;
thread_status[1024] = `IFUPATH256.swl.thr0_state;
thread_status[1025] = `IFUPATH256.swl.thr1_state;
thread_status[1026] = `IFUPATH256.swl.thr2_state;
thread_status[1027] = `IFUPATH256.swl.thr3_state;
thread_status[1028] = `IFUPATH257.swl.thr0_state;
thread_status[1029] = `IFUPATH257.swl.thr1_state;
thread_status[1030] = `IFUPATH257.swl.thr2_state;
thread_status[1031] = `IFUPATH257.swl.thr3_state;
thread_status[1032] = `IFUPATH258.swl.thr0_state;
thread_status[1033] = `IFUPATH258.swl.thr1_state;
thread_status[1034] = `IFUPATH258.swl.thr2_state;
thread_status[1035] = `IFUPATH258.swl.thr3_state;
thread_status[1036] = `IFUPATH259.swl.thr0_state;
thread_status[1037] = `IFUPATH259.swl.thr1_state;
thread_status[1038] = `IFUPATH259.swl.thr2_state;
thread_status[1039] = `IFUPATH259.swl.thr3_state;
thread_status[1040] = `IFUPATH260.swl.thr0_state;
thread_status[1041] = `IFUPATH260.swl.thr1_state;
thread_status[1042] = `IFUPATH260.swl.thr2_state;
thread_status[1043] = `IFUPATH260.swl.thr3_state;
thread_status[1044] = `IFUPATH261.swl.thr0_state;
thread_status[1045] = `IFUPATH261.swl.thr1_state;
thread_status[1046] = `IFUPATH261.swl.thr2_state;
thread_status[1047] = `IFUPATH261.swl.thr3_state;
thread_status[1048] = `IFUPATH262.swl.thr0_state;
thread_status[1049] = `IFUPATH262.swl.thr1_state;
thread_status[1050] = `IFUPATH262.swl.thr2_state;
thread_status[1051] = `IFUPATH262.swl.thr3_state;
thread_status[1052] = `IFUPATH263.swl.thr0_state;
thread_status[1053] = `IFUPATH263.swl.thr1_state;
thread_status[1054] = `IFUPATH263.swl.thr2_state;
thread_status[1055] = `IFUPATH263.swl.thr3_state;
thread_status[1056] = `IFUPATH264.swl.thr0_state;
thread_status[1057] = `IFUPATH264.swl.thr1_state;
thread_status[1058] = `IFUPATH264.swl.thr2_state;
thread_status[1059] = `IFUPATH264.swl.thr3_state;
thread_status[1060] = `IFUPATH265.swl.thr0_state;
thread_status[1061] = `IFUPATH265.swl.thr1_state;
thread_status[1062] = `IFUPATH265.swl.thr2_state;
thread_status[1063] = `IFUPATH265.swl.thr3_state;
thread_status[1064] = `IFUPATH266.swl.thr0_state;
thread_status[1065] = `IFUPATH266.swl.thr1_state;
thread_status[1066] = `IFUPATH266.swl.thr2_state;
thread_status[1067] = `IFUPATH266.swl.thr3_state;
thread_status[1068] = `IFUPATH267.swl.thr0_state;
thread_status[1069] = `IFUPATH267.swl.thr1_state;
thread_status[1070] = `IFUPATH267.swl.thr2_state;
thread_status[1071] = `IFUPATH267.swl.thr3_state;
thread_status[1072] = `IFUPATH268.swl.thr0_state;
thread_status[1073] = `IFUPATH268.swl.thr1_state;
thread_status[1074] = `IFUPATH268.swl.thr2_state;
thread_status[1075] = `IFUPATH268.swl.thr3_state;
thread_status[1076] = `IFUPATH269.swl.thr0_state;
thread_status[1077] = `IFUPATH269.swl.thr1_state;
thread_status[1078] = `IFUPATH269.swl.thr2_state;
thread_status[1079] = `IFUPATH269.swl.thr3_state;
thread_status[1080] = `IFUPATH270.swl.thr0_state;
thread_status[1081] = `IFUPATH270.swl.thr1_state;
thread_status[1082] = `IFUPATH270.swl.thr2_state;
thread_status[1083] = `IFUPATH270.swl.thr3_state;
thread_status[1084] = `IFUPATH271.swl.thr0_state;
thread_status[1085] = `IFUPATH271.swl.thr1_state;
thread_status[1086] = `IFUPATH271.swl.thr2_state;
thread_status[1087] = `IFUPATH271.swl.thr3_state;
thread_status[1088] = `IFUPATH272.swl.thr0_state;
thread_status[1089] = `IFUPATH272.swl.thr1_state;
thread_status[1090] = `IFUPATH272.swl.thr2_state;
thread_status[1091] = `IFUPATH272.swl.thr3_state;
thread_status[1092] = `IFUPATH273.swl.thr0_state;
thread_status[1093] = `IFUPATH273.swl.thr1_state;
thread_status[1094] = `IFUPATH273.swl.thr2_state;
thread_status[1095] = `IFUPATH273.swl.thr3_state;
thread_status[1096] = `IFUPATH274.swl.thr0_state;
thread_status[1097] = `IFUPATH274.swl.thr1_state;
thread_status[1098] = `IFUPATH274.swl.thr2_state;
thread_status[1099] = `IFUPATH274.swl.thr3_state;
thread_status[1100] = `IFUPATH275.swl.thr0_state;
thread_status[1101] = `IFUPATH275.swl.thr1_state;
thread_status[1102] = `IFUPATH275.swl.thr2_state;
thread_status[1103] = `IFUPATH275.swl.thr3_state;
thread_status[1104] = `IFUPATH276.swl.thr0_state;
thread_status[1105] = `IFUPATH276.swl.thr1_state;
thread_status[1106] = `IFUPATH276.swl.thr2_state;
thread_status[1107] = `IFUPATH276.swl.thr3_state;
thread_status[1108] = `IFUPATH277.swl.thr0_state;
thread_status[1109] = `IFUPATH277.swl.thr1_state;
thread_status[1110] = `IFUPATH277.swl.thr2_state;
thread_status[1111] = `IFUPATH277.swl.thr3_state;
thread_status[1112] = `IFUPATH278.swl.thr0_state;
thread_status[1113] = `IFUPATH278.swl.thr1_state;
thread_status[1114] = `IFUPATH278.swl.thr2_state;
thread_status[1115] = `IFUPATH278.swl.thr3_state;
thread_status[1116] = `IFUPATH279.swl.thr0_state;
thread_status[1117] = `IFUPATH279.swl.thr1_state;
thread_status[1118] = `IFUPATH279.swl.thr2_state;
thread_status[1119] = `IFUPATH279.swl.thr3_state;
thread_status[1120] = `IFUPATH280.swl.thr0_state;
thread_status[1121] = `IFUPATH280.swl.thr1_state;
thread_status[1122] = `IFUPATH280.swl.thr2_state;
thread_status[1123] = `IFUPATH280.swl.thr3_state;
thread_status[1124] = `IFUPATH281.swl.thr0_state;
thread_status[1125] = `IFUPATH281.swl.thr1_state;
thread_status[1126] = `IFUPATH281.swl.thr2_state;
thread_status[1127] = `IFUPATH281.swl.thr3_state;
thread_status[1128] = `IFUPATH282.swl.thr0_state;
thread_status[1129] = `IFUPATH282.swl.thr1_state;
thread_status[1130] = `IFUPATH282.swl.thr2_state;
thread_status[1131] = `IFUPATH282.swl.thr3_state;
thread_status[1132] = `IFUPATH283.swl.thr0_state;
thread_status[1133] = `IFUPATH283.swl.thr1_state;
thread_status[1134] = `IFUPATH283.swl.thr2_state;
thread_status[1135] = `IFUPATH283.swl.thr3_state;
thread_status[1136] = `IFUPATH284.swl.thr0_state;
thread_status[1137] = `IFUPATH284.swl.thr1_state;
thread_status[1138] = `IFUPATH284.swl.thr2_state;
thread_status[1139] = `IFUPATH284.swl.thr3_state;
thread_status[1140] = `IFUPATH285.swl.thr0_state;
thread_status[1141] = `IFUPATH285.swl.thr1_state;
thread_status[1142] = `IFUPATH285.swl.thr2_state;
thread_status[1143] = `IFUPATH285.swl.thr3_state;
thread_status[1144] = `IFUPATH286.swl.thr0_state;
thread_status[1145] = `IFUPATH286.swl.thr1_state;
thread_status[1146] = `IFUPATH286.swl.thr2_state;
thread_status[1147] = `IFUPATH286.swl.thr3_state;
thread_status[1148] = `IFUPATH287.swl.thr0_state;
thread_status[1149] = `IFUPATH287.swl.thr1_state;
thread_status[1150] = `IFUPATH287.swl.thr2_state;
thread_status[1151] = `IFUPATH287.swl.thr3_state;
thread_status[1152] = `IFUPATH288.swl.thr0_state;
thread_status[1153] = `IFUPATH288.swl.thr1_state;
thread_status[1154] = `IFUPATH288.swl.thr2_state;
thread_status[1155] = `IFUPATH288.swl.thr3_state;
thread_status[1156] = `IFUPATH289.swl.thr0_state;
thread_status[1157] = `IFUPATH289.swl.thr1_state;
thread_status[1158] = `IFUPATH289.swl.thr2_state;
thread_status[1159] = `IFUPATH289.swl.thr3_state;
thread_status[1160] = `IFUPATH290.swl.thr0_state;
thread_status[1161] = `IFUPATH290.swl.thr1_state;
thread_status[1162] = `IFUPATH290.swl.thr2_state;
thread_status[1163] = `IFUPATH290.swl.thr3_state;
thread_status[1164] = `IFUPATH291.swl.thr0_state;
thread_status[1165] = `IFUPATH291.swl.thr1_state;
thread_status[1166] = `IFUPATH291.swl.thr2_state;
thread_status[1167] = `IFUPATH291.swl.thr3_state;
thread_status[1168] = `IFUPATH292.swl.thr0_state;
thread_status[1169] = `IFUPATH292.swl.thr1_state;
thread_status[1170] = `IFUPATH292.swl.thr2_state;
thread_status[1171] = `IFUPATH292.swl.thr3_state;
thread_status[1172] = `IFUPATH293.swl.thr0_state;
thread_status[1173] = `IFUPATH293.swl.thr1_state;
thread_status[1174] = `IFUPATH293.swl.thr2_state;
thread_status[1175] = `IFUPATH293.swl.thr3_state;
thread_status[1176] = `IFUPATH294.swl.thr0_state;
thread_status[1177] = `IFUPATH294.swl.thr1_state;
thread_status[1178] = `IFUPATH294.swl.thr2_state;
thread_status[1179] = `IFUPATH294.swl.thr3_state;
thread_status[1180] = `IFUPATH295.swl.thr0_state;
thread_status[1181] = `IFUPATH295.swl.thr1_state;
thread_status[1182] = `IFUPATH295.swl.thr2_state;
thread_status[1183] = `IFUPATH295.swl.thr3_state;
thread_status[1184] = `IFUPATH296.swl.thr0_state;
thread_status[1185] = `IFUPATH296.swl.thr1_state;
thread_status[1186] = `IFUPATH296.swl.thr2_state;
thread_status[1187] = `IFUPATH296.swl.thr3_state;
thread_status[1188] = `IFUPATH297.swl.thr0_state;
thread_status[1189] = `IFUPATH297.swl.thr1_state;
thread_status[1190] = `IFUPATH297.swl.thr2_state;
thread_status[1191] = `IFUPATH297.swl.thr3_state;
thread_status[1192] = `IFUPATH298.swl.thr0_state;
thread_status[1193] = `IFUPATH298.swl.thr1_state;
thread_status[1194] = `IFUPATH298.swl.thr2_state;
thread_status[1195] = `IFUPATH298.swl.thr3_state;
thread_status[1196] = `IFUPATH299.swl.thr0_state;
thread_status[1197] = `IFUPATH299.swl.thr1_state;
thread_status[1198] = `IFUPATH299.swl.thr2_state;
thread_status[1199] = `IFUPATH299.swl.thr3_state;
thread_status[1200] = `IFUPATH300.swl.thr0_state;
thread_status[1201] = `IFUPATH300.swl.thr1_state;
thread_status[1202] = `IFUPATH300.swl.thr2_state;
thread_status[1203] = `IFUPATH300.swl.thr3_state;
thread_status[1204] = `IFUPATH301.swl.thr0_state;
thread_status[1205] = `IFUPATH301.swl.thr1_state;
thread_status[1206] = `IFUPATH301.swl.thr2_state;
thread_status[1207] = `IFUPATH301.swl.thr3_state;
thread_status[1208] = `IFUPATH302.swl.thr0_state;
thread_status[1209] = `IFUPATH302.swl.thr1_state;
thread_status[1210] = `IFUPATH302.swl.thr2_state;
thread_status[1211] = `IFUPATH302.swl.thr3_state;
thread_status[1212] = `IFUPATH303.swl.thr0_state;
thread_status[1213] = `IFUPATH303.swl.thr1_state;
thread_status[1214] = `IFUPATH303.swl.thr2_state;
thread_status[1215] = `IFUPATH303.swl.thr3_state;
thread_status[1216] = `IFUPATH304.swl.thr0_state;
thread_status[1217] = `IFUPATH304.swl.thr1_state;
thread_status[1218] = `IFUPATH304.swl.thr2_state;
thread_status[1219] = `IFUPATH304.swl.thr3_state;
thread_status[1220] = `IFUPATH305.swl.thr0_state;
thread_status[1221] = `IFUPATH305.swl.thr1_state;
thread_status[1222] = `IFUPATH305.swl.thr2_state;
thread_status[1223] = `IFUPATH305.swl.thr3_state;
thread_status[1224] = `IFUPATH306.swl.thr0_state;
thread_status[1225] = `IFUPATH306.swl.thr1_state;
thread_status[1226] = `IFUPATH306.swl.thr2_state;
thread_status[1227] = `IFUPATH306.swl.thr3_state;
thread_status[1228] = `IFUPATH307.swl.thr0_state;
thread_status[1229] = `IFUPATH307.swl.thr1_state;
thread_status[1230] = `IFUPATH307.swl.thr2_state;
thread_status[1231] = `IFUPATH307.swl.thr3_state;
thread_status[1232] = `IFUPATH308.swl.thr0_state;
thread_status[1233] = `IFUPATH308.swl.thr1_state;
thread_status[1234] = `IFUPATH308.swl.thr2_state;
thread_status[1235] = `IFUPATH308.swl.thr3_state;
thread_status[1236] = `IFUPATH309.swl.thr0_state;
thread_status[1237] = `IFUPATH309.swl.thr1_state;
thread_status[1238] = `IFUPATH309.swl.thr2_state;
thread_status[1239] = `IFUPATH309.swl.thr3_state;
thread_status[1240] = `IFUPATH310.swl.thr0_state;
thread_status[1241] = `IFUPATH310.swl.thr1_state;
thread_status[1242] = `IFUPATH310.swl.thr2_state;
thread_status[1243] = `IFUPATH310.swl.thr3_state;
thread_status[1244] = `IFUPATH311.swl.thr0_state;
thread_status[1245] = `IFUPATH311.swl.thr1_state;
thread_status[1246] = `IFUPATH311.swl.thr2_state;
thread_status[1247] = `IFUPATH311.swl.thr3_state;
thread_status[1248] = `IFUPATH312.swl.thr0_state;
thread_status[1249] = `IFUPATH312.swl.thr1_state;
thread_status[1250] = `IFUPATH312.swl.thr2_state;
thread_status[1251] = `IFUPATH312.swl.thr3_state;
thread_status[1252] = `IFUPATH313.swl.thr0_state;
thread_status[1253] = `IFUPATH313.swl.thr1_state;
thread_status[1254] = `IFUPATH313.swl.thr2_state;
thread_status[1255] = `IFUPATH313.swl.thr3_state;
thread_status[1256] = `IFUPATH314.swl.thr0_state;
thread_status[1257] = `IFUPATH314.swl.thr1_state;
thread_status[1258] = `IFUPATH314.swl.thr2_state;
thread_status[1259] = `IFUPATH314.swl.thr3_state;
thread_status[1260] = `IFUPATH315.swl.thr0_state;
thread_status[1261] = `IFUPATH315.swl.thr1_state;
thread_status[1262] = `IFUPATH315.swl.thr2_state;
thread_status[1263] = `IFUPATH315.swl.thr3_state;
thread_status[1264] = `IFUPATH316.swl.thr0_state;
thread_status[1265] = `IFUPATH316.swl.thr1_state;
thread_status[1266] = `IFUPATH316.swl.thr2_state;
thread_status[1267] = `IFUPATH316.swl.thr3_state;
thread_status[1268] = `IFUPATH317.swl.thr0_state;
thread_status[1269] = `IFUPATH317.swl.thr1_state;
thread_status[1270] = `IFUPATH317.swl.thr2_state;
thread_status[1271] = `IFUPATH317.swl.thr3_state;
thread_status[1272] = `IFUPATH318.swl.thr0_state;
thread_status[1273] = `IFUPATH318.swl.thr1_state;
thread_status[1274] = `IFUPATH318.swl.thr2_state;
thread_status[1275] = `IFUPATH318.swl.thr3_state;
thread_status[1276] = `IFUPATH319.swl.thr0_state;
thread_status[1277] = `IFUPATH319.swl.thr1_state;
thread_status[1278] = `IFUPATH319.swl.thr2_state;
thread_status[1279] = `IFUPATH319.swl.thr3_state;
thread_status[1280] = `IFUPATH320.swl.thr0_state;
thread_status[1281] = `IFUPATH320.swl.thr1_state;
thread_status[1282] = `IFUPATH320.swl.thr2_state;
thread_status[1283] = `IFUPATH320.swl.thr3_state;
thread_status[1284] = `IFUPATH321.swl.thr0_state;
thread_status[1285] = `IFUPATH321.swl.thr1_state;
thread_status[1286] = `IFUPATH321.swl.thr2_state;
thread_status[1287] = `IFUPATH321.swl.thr3_state;
thread_status[1288] = `IFUPATH322.swl.thr0_state;
thread_status[1289] = `IFUPATH322.swl.thr1_state;
thread_status[1290] = `IFUPATH322.swl.thr2_state;
thread_status[1291] = `IFUPATH322.swl.thr3_state;
thread_status[1292] = `IFUPATH323.swl.thr0_state;
thread_status[1293] = `IFUPATH323.swl.thr1_state;
thread_status[1294] = `IFUPATH323.swl.thr2_state;
thread_status[1295] = `IFUPATH323.swl.thr3_state;
thread_status[1296] = `IFUPATH324.swl.thr0_state;
thread_status[1297] = `IFUPATH324.swl.thr1_state;
thread_status[1298] = `IFUPATH324.swl.thr2_state;
thread_status[1299] = `IFUPATH324.swl.thr3_state;
thread_status[1300] = `IFUPATH325.swl.thr0_state;
thread_status[1301] = `IFUPATH325.swl.thr1_state;
thread_status[1302] = `IFUPATH325.swl.thr2_state;
thread_status[1303] = `IFUPATH325.swl.thr3_state;
thread_status[1304] = `IFUPATH326.swl.thr0_state;
thread_status[1305] = `IFUPATH326.swl.thr1_state;
thread_status[1306] = `IFUPATH326.swl.thr2_state;
thread_status[1307] = `IFUPATH326.swl.thr3_state;
thread_status[1308] = `IFUPATH327.swl.thr0_state;
thread_status[1309] = `IFUPATH327.swl.thr1_state;
thread_status[1310] = `IFUPATH327.swl.thr2_state;
thread_status[1311] = `IFUPATH327.swl.thr3_state;
thread_status[1312] = `IFUPATH328.swl.thr0_state;
thread_status[1313] = `IFUPATH328.swl.thr1_state;
thread_status[1314] = `IFUPATH328.swl.thr2_state;
thread_status[1315] = `IFUPATH328.swl.thr3_state;
thread_status[1316] = `IFUPATH329.swl.thr0_state;
thread_status[1317] = `IFUPATH329.swl.thr1_state;
thread_status[1318] = `IFUPATH329.swl.thr2_state;
thread_status[1319] = `IFUPATH329.swl.thr3_state;
thread_status[1320] = `IFUPATH330.swl.thr0_state;
thread_status[1321] = `IFUPATH330.swl.thr1_state;
thread_status[1322] = `IFUPATH330.swl.thr2_state;
thread_status[1323] = `IFUPATH330.swl.thr3_state;
thread_status[1324] = `IFUPATH331.swl.thr0_state;
thread_status[1325] = `IFUPATH331.swl.thr1_state;
thread_status[1326] = `IFUPATH331.swl.thr2_state;
thread_status[1327] = `IFUPATH331.swl.thr3_state;
thread_status[1328] = `IFUPATH332.swl.thr0_state;
thread_status[1329] = `IFUPATH332.swl.thr1_state;
thread_status[1330] = `IFUPATH332.swl.thr2_state;
thread_status[1331] = `IFUPATH332.swl.thr3_state;
thread_status[1332] = `IFUPATH333.swl.thr0_state;
thread_status[1333] = `IFUPATH333.swl.thr1_state;
thread_status[1334] = `IFUPATH333.swl.thr2_state;
thread_status[1335] = `IFUPATH333.swl.thr3_state;
thread_status[1336] = `IFUPATH334.swl.thr0_state;
thread_status[1337] = `IFUPATH334.swl.thr1_state;
thread_status[1338] = `IFUPATH334.swl.thr2_state;
thread_status[1339] = `IFUPATH334.swl.thr3_state;
thread_status[1340] = `IFUPATH335.swl.thr0_state;
thread_status[1341] = `IFUPATH335.swl.thr1_state;
thread_status[1342] = `IFUPATH335.swl.thr2_state;
thread_status[1343] = `IFUPATH335.swl.thr3_state;
thread_status[1344] = `IFUPATH336.swl.thr0_state;
thread_status[1345] = `IFUPATH336.swl.thr1_state;
thread_status[1346] = `IFUPATH336.swl.thr2_state;
thread_status[1347] = `IFUPATH336.swl.thr3_state;
thread_status[1348] = `IFUPATH337.swl.thr0_state;
thread_status[1349] = `IFUPATH337.swl.thr1_state;
thread_status[1350] = `IFUPATH337.swl.thr2_state;
thread_status[1351] = `IFUPATH337.swl.thr3_state;
thread_status[1352] = `IFUPATH338.swl.thr0_state;
thread_status[1353] = `IFUPATH338.swl.thr1_state;
thread_status[1354] = `IFUPATH338.swl.thr2_state;
thread_status[1355] = `IFUPATH338.swl.thr3_state;
thread_status[1356] = `IFUPATH339.swl.thr0_state;
thread_status[1357] = `IFUPATH339.swl.thr1_state;
thread_status[1358] = `IFUPATH339.swl.thr2_state;
thread_status[1359] = `IFUPATH339.swl.thr3_state;
thread_status[1360] = `IFUPATH340.swl.thr0_state;
thread_status[1361] = `IFUPATH340.swl.thr1_state;
thread_status[1362] = `IFUPATH340.swl.thr2_state;
thread_status[1363] = `IFUPATH340.swl.thr3_state;
thread_status[1364] = `IFUPATH341.swl.thr0_state;
thread_status[1365] = `IFUPATH341.swl.thr1_state;
thread_status[1366] = `IFUPATH341.swl.thr2_state;
thread_status[1367] = `IFUPATH341.swl.thr3_state;
thread_status[1368] = `IFUPATH342.swl.thr0_state;
thread_status[1369] = `IFUPATH342.swl.thr1_state;
thread_status[1370] = `IFUPATH342.swl.thr2_state;
thread_status[1371] = `IFUPATH342.swl.thr3_state;
thread_status[1372] = `IFUPATH343.swl.thr0_state;
thread_status[1373] = `IFUPATH343.swl.thr1_state;
thread_status[1374] = `IFUPATH343.swl.thr2_state;
thread_status[1375] = `IFUPATH343.swl.thr3_state;
thread_status[1376] = `IFUPATH344.swl.thr0_state;
thread_status[1377] = `IFUPATH344.swl.thr1_state;
thread_status[1378] = `IFUPATH344.swl.thr2_state;
thread_status[1379] = `IFUPATH344.swl.thr3_state;
thread_status[1380] = `IFUPATH345.swl.thr0_state;
thread_status[1381] = `IFUPATH345.swl.thr1_state;
thread_status[1382] = `IFUPATH345.swl.thr2_state;
thread_status[1383] = `IFUPATH345.swl.thr3_state;
thread_status[1384] = `IFUPATH346.swl.thr0_state;
thread_status[1385] = `IFUPATH346.swl.thr1_state;
thread_status[1386] = `IFUPATH346.swl.thr2_state;
thread_status[1387] = `IFUPATH346.swl.thr3_state;
thread_status[1388] = `IFUPATH347.swl.thr0_state;
thread_status[1389] = `IFUPATH347.swl.thr1_state;
thread_status[1390] = `IFUPATH347.swl.thr2_state;
thread_status[1391] = `IFUPATH347.swl.thr3_state;
thread_status[1392] = `IFUPATH348.swl.thr0_state;
thread_status[1393] = `IFUPATH348.swl.thr1_state;
thread_status[1394] = `IFUPATH348.swl.thr2_state;
thread_status[1395] = `IFUPATH348.swl.thr3_state;
thread_status[1396] = `IFUPATH349.swl.thr0_state;
thread_status[1397] = `IFUPATH349.swl.thr1_state;
thread_status[1398] = `IFUPATH349.swl.thr2_state;
thread_status[1399] = `IFUPATH349.swl.thr3_state;
thread_status[1400] = `IFUPATH350.swl.thr0_state;
thread_status[1401] = `IFUPATH350.swl.thr1_state;
thread_status[1402] = `IFUPATH350.swl.thr2_state;
thread_status[1403] = `IFUPATH350.swl.thr3_state;
thread_status[1404] = `IFUPATH351.swl.thr0_state;
thread_status[1405] = `IFUPATH351.swl.thr1_state;
thread_status[1406] = `IFUPATH351.swl.thr2_state;
thread_status[1407] = `IFUPATH351.swl.thr3_state;
thread_status[1408] = `IFUPATH352.swl.thr0_state;
thread_status[1409] = `IFUPATH352.swl.thr1_state;
thread_status[1410] = `IFUPATH352.swl.thr2_state;
thread_status[1411] = `IFUPATH352.swl.thr3_state;
thread_status[1412] = `IFUPATH353.swl.thr0_state;
thread_status[1413] = `IFUPATH353.swl.thr1_state;
thread_status[1414] = `IFUPATH353.swl.thr2_state;
thread_status[1415] = `IFUPATH353.swl.thr3_state;
thread_status[1416] = `IFUPATH354.swl.thr0_state;
thread_status[1417] = `IFUPATH354.swl.thr1_state;
thread_status[1418] = `IFUPATH354.swl.thr2_state;
thread_status[1419] = `IFUPATH354.swl.thr3_state;
thread_status[1420] = `IFUPATH355.swl.thr0_state;
thread_status[1421] = `IFUPATH355.swl.thr1_state;
thread_status[1422] = `IFUPATH355.swl.thr2_state;
thread_status[1423] = `IFUPATH355.swl.thr3_state;
thread_status[1424] = `IFUPATH356.swl.thr0_state;
thread_status[1425] = `IFUPATH356.swl.thr1_state;
thread_status[1426] = `IFUPATH356.swl.thr2_state;
thread_status[1427] = `IFUPATH356.swl.thr3_state;
thread_status[1428] = `IFUPATH357.swl.thr0_state;
thread_status[1429] = `IFUPATH357.swl.thr1_state;
thread_status[1430] = `IFUPATH357.swl.thr2_state;
thread_status[1431] = `IFUPATH357.swl.thr3_state;
thread_status[1432] = `IFUPATH358.swl.thr0_state;
thread_status[1433] = `IFUPATH358.swl.thr1_state;
thread_status[1434] = `IFUPATH358.swl.thr2_state;
thread_status[1435] = `IFUPATH358.swl.thr3_state;
thread_status[1436] = `IFUPATH359.swl.thr0_state;
thread_status[1437] = `IFUPATH359.swl.thr1_state;
thread_status[1438] = `IFUPATH359.swl.thr2_state;
thread_status[1439] = `IFUPATH359.swl.thr3_state;
thread_status[1440] = `IFUPATH360.swl.thr0_state;
thread_status[1441] = `IFUPATH360.swl.thr1_state;
thread_status[1442] = `IFUPATH360.swl.thr2_state;
thread_status[1443] = `IFUPATH360.swl.thr3_state;
thread_status[1444] = `IFUPATH361.swl.thr0_state;
thread_status[1445] = `IFUPATH361.swl.thr1_state;
thread_status[1446] = `IFUPATH361.swl.thr2_state;
thread_status[1447] = `IFUPATH361.swl.thr3_state;
thread_status[1448] = `IFUPATH362.swl.thr0_state;
thread_status[1449] = `IFUPATH362.swl.thr1_state;
thread_status[1450] = `IFUPATH362.swl.thr2_state;
thread_status[1451] = `IFUPATH362.swl.thr3_state;
thread_status[1452] = `IFUPATH363.swl.thr0_state;
thread_status[1453] = `IFUPATH363.swl.thr1_state;
thread_status[1454] = `IFUPATH363.swl.thr2_state;
thread_status[1455] = `IFUPATH363.swl.thr3_state;
thread_status[1456] = `IFUPATH364.swl.thr0_state;
thread_status[1457] = `IFUPATH364.swl.thr1_state;
thread_status[1458] = `IFUPATH364.swl.thr2_state;
thread_status[1459] = `IFUPATH364.swl.thr3_state;
thread_status[1460] = `IFUPATH365.swl.thr0_state;
thread_status[1461] = `IFUPATH365.swl.thr1_state;
thread_status[1462] = `IFUPATH365.swl.thr2_state;
thread_status[1463] = `IFUPATH365.swl.thr3_state;
thread_status[1464] = `IFUPATH366.swl.thr0_state;
thread_status[1465] = `IFUPATH366.swl.thr1_state;
thread_status[1466] = `IFUPATH366.swl.thr2_state;
thread_status[1467] = `IFUPATH366.swl.thr3_state;
thread_status[1468] = `IFUPATH367.swl.thr0_state;
thread_status[1469] = `IFUPATH367.swl.thr1_state;
thread_status[1470] = `IFUPATH367.swl.thr2_state;
thread_status[1471] = `IFUPATH367.swl.thr3_state;
thread_status[1472] = `IFUPATH368.swl.thr0_state;
thread_status[1473] = `IFUPATH368.swl.thr1_state;
thread_status[1474] = `IFUPATH368.swl.thr2_state;
thread_status[1475] = `IFUPATH368.swl.thr3_state;
thread_status[1476] = `IFUPATH369.swl.thr0_state;
thread_status[1477] = `IFUPATH369.swl.thr1_state;
thread_status[1478] = `IFUPATH369.swl.thr2_state;
thread_status[1479] = `IFUPATH369.swl.thr3_state;
thread_status[1480] = `IFUPATH370.swl.thr0_state;
thread_status[1481] = `IFUPATH370.swl.thr1_state;
thread_status[1482] = `IFUPATH370.swl.thr2_state;
thread_status[1483] = `IFUPATH370.swl.thr3_state;
thread_status[1484] = `IFUPATH371.swl.thr0_state;
thread_status[1485] = `IFUPATH371.swl.thr1_state;
thread_status[1486] = `IFUPATH371.swl.thr2_state;
thread_status[1487] = `IFUPATH371.swl.thr3_state;
thread_status[1488] = `IFUPATH372.swl.thr0_state;
thread_status[1489] = `IFUPATH372.swl.thr1_state;
thread_status[1490] = `IFUPATH372.swl.thr2_state;
thread_status[1491] = `IFUPATH372.swl.thr3_state;
thread_status[1492] = `IFUPATH373.swl.thr0_state;
thread_status[1493] = `IFUPATH373.swl.thr1_state;
thread_status[1494] = `IFUPATH373.swl.thr2_state;
thread_status[1495] = `IFUPATH373.swl.thr3_state;
thread_status[1496] = `IFUPATH374.swl.thr0_state;
thread_status[1497] = `IFUPATH374.swl.thr1_state;
thread_status[1498] = `IFUPATH374.swl.thr2_state;
thread_status[1499] = `IFUPATH374.swl.thr3_state;
thread_status[1500] = `IFUPATH375.swl.thr0_state;
thread_status[1501] = `IFUPATH375.swl.thr1_state;
thread_status[1502] = `IFUPATH375.swl.thr2_state;
thread_status[1503] = `IFUPATH375.swl.thr3_state;
thread_status[1504] = `IFUPATH376.swl.thr0_state;
thread_status[1505] = `IFUPATH376.swl.thr1_state;
thread_status[1506] = `IFUPATH376.swl.thr2_state;
thread_status[1507] = `IFUPATH376.swl.thr3_state;
thread_status[1508] = `IFUPATH377.swl.thr0_state;
thread_status[1509] = `IFUPATH377.swl.thr1_state;
thread_status[1510] = `IFUPATH377.swl.thr2_state;
thread_status[1511] = `IFUPATH377.swl.thr3_state;
thread_status[1512] = `IFUPATH378.swl.thr0_state;
thread_status[1513] = `IFUPATH378.swl.thr1_state;
thread_status[1514] = `IFUPATH378.swl.thr2_state;
thread_status[1515] = `IFUPATH378.swl.thr3_state;
thread_status[1516] = `IFUPATH379.swl.thr0_state;
thread_status[1517] = `IFUPATH379.swl.thr1_state;
thread_status[1518] = `IFUPATH379.swl.thr2_state;
thread_status[1519] = `IFUPATH379.swl.thr3_state;
thread_status[1520] = `IFUPATH380.swl.thr0_state;
thread_status[1521] = `IFUPATH380.swl.thr1_state;
thread_status[1522] = `IFUPATH380.swl.thr2_state;
thread_status[1523] = `IFUPATH380.swl.thr3_state;
thread_status[1524] = `IFUPATH381.swl.thr0_state;
thread_status[1525] = `IFUPATH381.swl.thr1_state;
thread_status[1526] = `IFUPATH381.swl.thr2_state;
thread_status[1527] = `IFUPATH381.swl.thr3_state;
thread_status[1528] = `IFUPATH382.swl.thr0_state;
thread_status[1529] = `IFUPATH382.swl.thr1_state;
thread_status[1530] = `IFUPATH382.swl.thr2_state;
thread_status[1531] = `IFUPATH382.swl.thr3_state;
thread_status[1532] = `IFUPATH383.swl.thr0_state;
thread_status[1533] = `IFUPATH383.swl.thr1_state;
thread_status[1534] = `IFUPATH383.swl.thr2_state;
thread_status[1535] = `IFUPATH383.swl.thr3_state;
thread_status[1536] = `IFUPATH384.swl.thr0_state;
thread_status[1537] = `IFUPATH384.swl.thr1_state;
thread_status[1538] = `IFUPATH384.swl.thr2_state;
thread_status[1539] = `IFUPATH384.swl.thr3_state;
thread_status[1540] = `IFUPATH385.swl.thr0_state;
thread_status[1541] = `IFUPATH385.swl.thr1_state;
thread_status[1542] = `IFUPATH385.swl.thr2_state;
thread_status[1543] = `IFUPATH385.swl.thr3_state;
thread_status[1544] = `IFUPATH386.swl.thr0_state;
thread_status[1545] = `IFUPATH386.swl.thr1_state;
thread_status[1546] = `IFUPATH386.swl.thr2_state;
thread_status[1547] = `IFUPATH386.swl.thr3_state;
thread_status[1548] = `IFUPATH387.swl.thr0_state;
thread_status[1549] = `IFUPATH387.swl.thr1_state;
thread_status[1550] = `IFUPATH387.swl.thr2_state;
thread_status[1551] = `IFUPATH387.swl.thr3_state;
thread_status[1552] = `IFUPATH388.swl.thr0_state;
thread_status[1553] = `IFUPATH388.swl.thr1_state;
thread_status[1554] = `IFUPATH388.swl.thr2_state;
thread_status[1555] = `IFUPATH388.swl.thr3_state;
thread_status[1556] = `IFUPATH389.swl.thr0_state;
thread_status[1557] = `IFUPATH389.swl.thr1_state;
thread_status[1558] = `IFUPATH389.swl.thr2_state;
thread_status[1559] = `IFUPATH389.swl.thr3_state;
thread_status[1560] = `IFUPATH390.swl.thr0_state;
thread_status[1561] = `IFUPATH390.swl.thr1_state;
thread_status[1562] = `IFUPATH390.swl.thr2_state;
thread_status[1563] = `IFUPATH390.swl.thr3_state;
thread_status[1564] = `IFUPATH391.swl.thr0_state;
thread_status[1565] = `IFUPATH391.swl.thr1_state;
thread_status[1566] = `IFUPATH391.swl.thr2_state;
thread_status[1567] = `IFUPATH391.swl.thr3_state;
thread_status[1568] = `IFUPATH392.swl.thr0_state;
thread_status[1569] = `IFUPATH392.swl.thr1_state;
thread_status[1570] = `IFUPATH392.swl.thr2_state;
thread_status[1571] = `IFUPATH392.swl.thr3_state;
thread_status[1572] = `IFUPATH393.swl.thr0_state;
thread_status[1573] = `IFUPATH393.swl.thr1_state;
thread_status[1574] = `IFUPATH393.swl.thr2_state;
thread_status[1575] = `IFUPATH393.swl.thr3_state;
thread_status[1576] = `IFUPATH394.swl.thr0_state;
thread_status[1577] = `IFUPATH394.swl.thr1_state;
thread_status[1578] = `IFUPATH394.swl.thr2_state;
thread_status[1579] = `IFUPATH394.swl.thr3_state;
thread_status[1580] = `IFUPATH395.swl.thr0_state;
thread_status[1581] = `IFUPATH395.swl.thr1_state;
thread_status[1582] = `IFUPATH395.swl.thr2_state;
thread_status[1583] = `IFUPATH395.swl.thr3_state;
thread_status[1584] = `IFUPATH396.swl.thr0_state;
thread_status[1585] = `IFUPATH396.swl.thr1_state;
thread_status[1586] = `IFUPATH396.swl.thr2_state;
thread_status[1587] = `IFUPATH396.swl.thr3_state;
thread_status[1588] = `IFUPATH397.swl.thr0_state;
thread_status[1589] = `IFUPATH397.swl.thr1_state;
thread_status[1590] = `IFUPATH397.swl.thr2_state;
thread_status[1591] = `IFUPATH397.swl.thr3_state;
thread_status[1592] = `IFUPATH398.swl.thr0_state;
thread_status[1593] = `IFUPATH398.swl.thr1_state;
thread_status[1594] = `IFUPATH398.swl.thr2_state;
thread_status[1595] = `IFUPATH398.swl.thr3_state;
thread_status[1596] = `IFUPATH399.swl.thr0_state;
thread_status[1597] = `IFUPATH399.swl.thr1_state;
thread_status[1598] = `IFUPATH399.swl.thr2_state;
thread_status[1599] = `IFUPATH399.swl.thr3_state;
thread_status[1600] = `IFUPATH400.swl.thr0_state;
thread_status[1601] = `IFUPATH400.swl.thr1_state;
thread_status[1602] = `IFUPATH400.swl.thr2_state;
thread_status[1603] = `IFUPATH400.swl.thr3_state;
thread_status[1604] = `IFUPATH401.swl.thr0_state;
thread_status[1605] = `IFUPATH401.swl.thr1_state;
thread_status[1606] = `IFUPATH401.swl.thr2_state;
thread_status[1607] = `IFUPATH401.swl.thr3_state;
thread_status[1608] = `IFUPATH402.swl.thr0_state;
thread_status[1609] = `IFUPATH402.swl.thr1_state;
thread_status[1610] = `IFUPATH402.swl.thr2_state;
thread_status[1611] = `IFUPATH402.swl.thr3_state;
thread_status[1612] = `IFUPATH403.swl.thr0_state;
thread_status[1613] = `IFUPATH403.swl.thr1_state;
thread_status[1614] = `IFUPATH403.swl.thr2_state;
thread_status[1615] = `IFUPATH403.swl.thr3_state;
thread_status[1616] = `IFUPATH404.swl.thr0_state;
thread_status[1617] = `IFUPATH404.swl.thr1_state;
thread_status[1618] = `IFUPATH404.swl.thr2_state;
thread_status[1619] = `IFUPATH404.swl.thr3_state;
thread_status[1620] = `IFUPATH405.swl.thr0_state;
thread_status[1621] = `IFUPATH405.swl.thr1_state;
thread_status[1622] = `IFUPATH405.swl.thr2_state;
thread_status[1623] = `IFUPATH405.swl.thr3_state;
thread_status[1624] = `IFUPATH406.swl.thr0_state;
thread_status[1625] = `IFUPATH406.swl.thr1_state;
thread_status[1626] = `IFUPATH406.swl.thr2_state;
thread_status[1627] = `IFUPATH406.swl.thr3_state;
thread_status[1628] = `IFUPATH407.swl.thr0_state;
thread_status[1629] = `IFUPATH407.swl.thr1_state;
thread_status[1630] = `IFUPATH407.swl.thr2_state;
thread_status[1631] = `IFUPATH407.swl.thr3_state;
thread_status[1632] = `IFUPATH408.swl.thr0_state;
thread_status[1633] = `IFUPATH408.swl.thr1_state;
thread_status[1634] = `IFUPATH408.swl.thr2_state;
thread_status[1635] = `IFUPATH408.swl.thr3_state;
thread_status[1636] = `IFUPATH409.swl.thr0_state;
thread_status[1637] = `IFUPATH409.swl.thr1_state;
thread_status[1638] = `IFUPATH409.swl.thr2_state;
thread_status[1639] = `IFUPATH409.swl.thr3_state;
thread_status[1640] = `IFUPATH410.swl.thr0_state;
thread_status[1641] = `IFUPATH410.swl.thr1_state;
thread_status[1642] = `IFUPATH410.swl.thr2_state;
thread_status[1643] = `IFUPATH410.swl.thr3_state;
thread_status[1644] = `IFUPATH411.swl.thr0_state;
thread_status[1645] = `IFUPATH411.swl.thr1_state;
thread_status[1646] = `IFUPATH411.swl.thr2_state;
thread_status[1647] = `IFUPATH411.swl.thr3_state;
thread_status[1648] = `IFUPATH412.swl.thr0_state;
thread_status[1649] = `IFUPATH412.swl.thr1_state;
thread_status[1650] = `IFUPATH412.swl.thr2_state;
thread_status[1651] = `IFUPATH412.swl.thr3_state;
thread_status[1652] = `IFUPATH413.swl.thr0_state;
thread_status[1653] = `IFUPATH413.swl.thr1_state;
thread_status[1654] = `IFUPATH413.swl.thr2_state;
thread_status[1655] = `IFUPATH413.swl.thr3_state;
thread_status[1656] = `IFUPATH414.swl.thr0_state;
thread_status[1657] = `IFUPATH414.swl.thr1_state;
thread_status[1658] = `IFUPATH414.swl.thr2_state;
thread_status[1659] = `IFUPATH414.swl.thr3_state;
thread_status[1660] = `IFUPATH415.swl.thr0_state;
thread_status[1661] = `IFUPATH415.swl.thr1_state;
thread_status[1662] = `IFUPATH415.swl.thr2_state;
thread_status[1663] = `IFUPATH415.swl.thr3_state;
thread_status[1664] = `IFUPATH416.swl.thr0_state;
thread_status[1665] = `IFUPATH416.swl.thr1_state;
thread_status[1666] = `IFUPATH416.swl.thr2_state;
thread_status[1667] = `IFUPATH416.swl.thr3_state;
thread_status[1668] = `IFUPATH417.swl.thr0_state;
thread_status[1669] = `IFUPATH417.swl.thr1_state;
thread_status[1670] = `IFUPATH417.swl.thr2_state;
thread_status[1671] = `IFUPATH417.swl.thr3_state;
thread_status[1672] = `IFUPATH418.swl.thr0_state;
thread_status[1673] = `IFUPATH418.swl.thr1_state;
thread_status[1674] = `IFUPATH418.swl.thr2_state;
thread_status[1675] = `IFUPATH418.swl.thr3_state;
thread_status[1676] = `IFUPATH419.swl.thr0_state;
thread_status[1677] = `IFUPATH419.swl.thr1_state;
thread_status[1678] = `IFUPATH419.swl.thr2_state;
thread_status[1679] = `IFUPATH419.swl.thr3_state;
thread_status[1680] = `IFUPATH420.swl.thr0_state;
thread_status[1681] = `IFUPATH420.swl.thr1_state;
thread_status[1682] = `IFUPATH420.swl.thr2_state;
thread_status[1683] = `IFUPATH420.swl.thr3_state;
thread_status[1684] = `IFUPATH421.swl.thr0_state;
thread_status[1685] = `IFUPATH421.swl.thr1_state;
thread_status[1686] = `IFUPATH421.swl.thr2_state;
thread_status[1687] = `IFUPATH421.swl.thr3_state;
thread_status[1688] = `IFUPATH422.swl.thr0_state;
thread_status[1689] = `IFUPATH422.swl.thr1_state;
thread_status[1690] = `IFUPATH422.swl.thr2_state;
thread_status[1691] = `IFUPATH422.swl.thr3_state;
thread_status[1692] = `IFUPATH423.swl.thr0_state;
thread_status[1693] = `IFUPATH423.swl.thr1_state;
thread_status[1694] = `IFUPATH423.swl.thr2_state;
thread_status[1695] = `IFUPATH423.swl.thr3_state;
thread_status[1696] = `IFUPATH424.swl.thr0_state;
thread_status[1697] = `IFUPATH424.swl.thr1_state;
thread_status[1698] = `IFUPATH424.swl.thr2_state;
thread_status[1699] = `IFUPATH424.swl.thr3_state;
thread_status[1700] = `IFUPATH425.swl.thr0_state;
thread_status[1701] = `IFUPATH425.swl.thr1_state;
thread_status[1702] = `IFUPATH425.swl.thr2_state;
thread_status[1703] = `IFUPATH425.swl.thr3_state;
thread_status[1704] = `IFUPATH426.swl.thr0_state;
thread_status[1705] = `IFUPATH426.swl.thr1_state;
thread_status[1706] = `IFUPATH426.swl.thr2_state;
thread_status[1707] = `IFUPATH426.swl.thr3_state;
thread_status[1708] = `IFUPATH427.swl.thr0_state;
thread_status[1709] = `IFUPATH427.swl.thr1_state;
thread_status[1710] = `IFUPATH427.swl.thr2_state;
thread_status[1711] = `IFUPATH427.swl.thr3_state;
thread_status[1712] = `IFUPATH428.swl.thr0_state;
thread_status[1713] = `IFUPATH428.swl.thr1_state;
thread_status[1714] = `IFUPATH428.swl.thr2_state;
thread_status[1715] = `IFUPATH428.swl.thr3_state;
thread_status[1716] = `IFUPATH429.swl.thr0_state;
thread_status[1717] = `IFUPATH429.swl.thr1_state;
thread_status[1718] = `IFUPATH429.swl.thr2_state;
thread_status[1719] = `IFUPATH429.swl.thr3_state;
thread_status[1720] = `IFUPATH430.swl.thr0_state;
thread_status[1721] = `IFUPATH430.swl.thr1_state;
thread_status[1722] = `IFUPATH430.swl.thr2_state;
thread_status[1723] = `IFUPATH430.swl.thr3_state;
thread_status[1724] = `IFUPATH431.swl.thr0_state;
thread_status[1725] = `IFUPATH431.swl.thr1_state;
thread_status[1726] = `IFUPATH431.swl.thr2_state;
thread_status[1727] = `IFUPATH431.swl.thr3_state;
thread_status[1728] = `IFUPATH432.swl.thr0_state;
thread_status[1729] = `IFUPATH432.swl.thr1_state;
thread_status[1730] = `IFUPATH432.swl.thr2_state;
thread_status[1731] = `IFUPATH432.swl.thr3_state;
thread_status[1732] = `IFUPATH433.swl.thr0_state;
thread_status[1733] = `IFUPATH433.swl.thr1_state;
thread_status[1734] = `IFUPATH433.swl.thr2_state;
thread_status[1735] = `IFUPATH433.swl.thr3_state;
thread_status[1736] = `IFUPATH434.swl.thr0_state;
thread_status[1737] = `IFUPATH434.swl.thr1_state;
thread_status[1738] = `IFUPATH434.swl.thr2_state;
thread_status[1739] = `IFUPATH434.swl.thr3_state;
thread_status[1740] = `IFUPATH435.swl.thr0_state;
thread_status[1741] = `IFUPATH435.swl.thr1_state;
thread_status[1742] = `IFUPATH435.swl.thr2_state;
thread_status[1743] = `IFUPATH435.swl.thr3_state;
thread_status[1744] = `IFUPATH436.swl.thr0_state;
thread_status[1745] = `IFUPATH436.swl.thr1_state;
thread_status[1746] = `IFUPATH436.swl.thr2_state;
thread_status[1747] = `IFUPATH436.swl.thr3_state;
thread_status[1748] = `IFUPATH437.swl.thr0_state;
thread_status[1749] = `IFUPATH437.swl.thr1_state;
thread_status[1750] = `IFUPATH437.swl.thr2_state;
thread_status[1751] = `IFUPATH437.swl.thr3_state;
thread_status[1752] = `IFUPATH438.swl.thr0_state;
thread_status[1753] = `IFUPATH438.swl.thr1_state;
thread_status[1754] = `IFUPATH438.swl.thr2_state;
thread_status[1755] = `IFUPATH438.swl.thr3_state;
thread_status[1756] = `IFUPATH439.swl.thr0_state;
thread_status[1757] = `IFUPATH439.swl.thr1_state;
thread_status[1758] = `IFUPATH439.swl.thr2_state;
thread_status[1759] = `IFUPATH439.swl.thr3_state;
thread_status[1760] = `IFUPATH440.swl.thr0_state;
thread_status[1761] = `IFUPATH440.swl.thr1_state;
thread_status[1762] = `IFUPATH440.swl.thr2_state;
thread_status[1763] = `IFUPATH440.swl.thr3_state;
thread_status[1764] = `IFUPATH441.swl.thr0_state;
thread_status[1765] = `IFUPATH441.swl.thr1_state;
thread_status[1766] = `IFUPATH441.swl.thr2_state;
thread_status[1767] = `IFUPATH441.swl.thr3_state;
thread_status[1768] = `IFUPATH442.swl.thr0_state;
thread_status[1769] = `IFUPATH442.swl.thr1_state;
thread_status[1770] = `IFUPATH442.swl.thr2_state;
thread_status[1771] = `IFUPATH442.swl.thr3_state;
thread_status[1772] = `IFUPATH443.swl.thr0_state;
thread_status[1773] = `IFUPATH443.swl.thr1_state;
thread_status[1774] = `IFUPATH443.swl.thr2_state;
thread_status[1775] = `IFUPATH443.swl.thr3_state;
thread_status[1776] = `IFUPATH444.swl.thr0_state;
thread_status[1777] = `IFUPATH444.swl.thr1_state;
thread_status[1778] = `IFUPATH444.swl.thr2_state;
thread_status[1779] = `IFUPATH444.swl.thr3_state;
thread_status[1780] = `IFUPATH445.swl.thr0_state;
thread_status[1781] = `IFUPATH445.swl.thr1_state;
thread_status[1782] = `IFUPATH445.swl.thr2_state;
thread_status[1783] = `IFUPATH445.swl.thr3_state;
thread_status[1784] = `IFUPATH446.swl.thr0_state;
thread_status[1785] = `IFUPATH446.swl.thr1_state;
thread_status[1786] = `IFUPATH446.swl.thr2_state;
thread_status[1787] = `IFUPATH446.swl.thr3_state;
thread_status[1788] = `IFUPATH447.swl.thr0_state;
thread_status[1789] = `IFUPATH447.swl.thr1_state;
thread_status[1790] = `IFUPATH447.swl.thr2_state;
thread_status[1791] = `IFUPATH447.swl.thr3_state;
thread_status[1792] = `IFUPATH448.swl.thr0_state;
thread_status[1793] = `IFUPATH448.swl.thr1_state;
thread_status[1794] = `IFUPATH448.swl.thr2_state;
thread_status[1795] = `IFUPATH448.swl.thr3_state;
thread_status[1796] = `IFUPATH449.swl.thr0_state;
thread_status[1797] = `IFUPATH449.swl.thr1_state;
thread_status[1798] = `IFUPATH449.swl.thr2_state;
thread_status[1799] = `IFUPATH449.swl.thr3_state;
thread_status[1800] = `IFUPATH450.swl.thr0_state;
thread_status[1801] = `IFUPATH450.swl.thr1_state;
thread_status[1802] = `IFUPATH450.swl.thr2_state;
thread_status[1803] = `IFUPATH450.swl.thr3_state;
thread_status[1804] = `IFUPATH451.swl.thr0_state;
thread_status[1805] = `IFUPATH451.swl.thr1_state;
thread_status[1806] = `IFUPATH451.swl.thr2_state;
thread_status[1807] = `IFUPATH451.swl.thr3_state;
thread_status[1808] = `IFUPATH452.swl.thr0_state;
thread_status[1809] = `IFUPATH452.swl.thr1_state;
thread_status[1810] = `IFUPATH452.swl.thr2_state;
thread_status[1811] = `IFUPATH452.swl.thr3_state;
thread_status[1812] = `IFUPATH453.swl.thr0_state;
thread_status[1813] = `IFUPATH453.swl.thr1_state;
thread_status[1814] = `IFUPATH453.swl.thr2_state;
thread_status[1815] = `IFUPATH453.swl.thr3_state;
thread_status[1816] = `IFUPATH454.swl.thr0_state;
thread_status[1817] = `IFUPATH454.swl.thr1_state;
thread_status[1818] = `IFUPATH454.swl.thr2_state;
thread_status[1819] = `IFUPATH454.swl.thr3_state;
thread_status[1820] = `IFUPATH455.swl.thr0_state;
thread_status[1821] = `IFUPATH455.swl.thr1_state;
thread_status[1822] = `IFUPATH455.swl.thr2_state;
thread_status[1823] = `IFUPATH455.swl.thr3_state;
thread_status[1824] = `IFUPATH456.swl.thr0_state;
thread_status[1825] = `IFUPATH456.swl.thr1_state;
thread_status[1826] = `IFUPATH456.swl.thr2_state;
thread_status[1827] = `IFUPATH456.swl.thr3_state;
thread_status[1828] = `IFUPATH457.swl.thr0_state;
thread_status[1829] = `IFUPATH457.swl.thr1_state;
thread_status[1830] = `IFUPATH457.swl.thr2_state;
thread_status[1831] = `IFUPATH457.swl.thr3_state;
thread_status[1832] = `IFUPATH458.swl.thr0_state;
thread_status[1833] = `IFUPATH458.swl.thr1_state;
thread_status[1834] = `IFUPATH458.swl.thr2_state;
thread_status[1835] = `IFUPATH458.swl.thr3_state;
thread_status[1836] = `IFUPATH459.swl.thr0_state;
thread_status[1837] = `IFUPATH459.swl.thr1_state;
thread_status[1838] = `IFUPATH459.swl.thr2_state;
thread_status[1839] = `IFUPATH459.swl.thr3_state;
thread_status[1840] = `IFUPATH460.swl.thr0_state;
thread_status[1841] = `IFUPATH460.swl.thr1_state;
thread_status[1842] = `IFUPATH460.swl.thr2_state;
thread_status[1843] = `IFUPATH460.swl.thr3_state;
thread_status[1844] = `IFUPATH461.swl.thr0_state;
thread_status[1845] = `IFUPATH461.swl.thr1_state;
thread_status[1846] = `IFUPATH461.swl.thr2_state;
thread_status[1847] = `IFUPATH461.swl.thr3_state;
thread_status[1848] = `IFUPATH462.swl.thr0_state;
thread_status[1849] = `IFUPATH462.swl.thr1_state;
thread_status[1850] = `IFUPATH462.swl.thr2_state;
thread_status[1851] = `IFUPATH462.swl.thr3_state;
thread_status[1852] = `IFUPATH463.swl.thr0_state;
thread_status[1853] = `IFUPATH463.swl.thr1_state;
thread_status[1854] = `IFUPATH463.swl.thr2_state;
thread_status[1855] = `IFUPATH463.swl.thr3_state;
thread_status[1856] = `IFUPATH464.swl.thr0_state;
thread_status[1857] = `IFUPATH464.swl.thr1_state;
thread_status[1858] = `IFUPATH464.swl.thr2_state;
thread_status[1859] = `IFUPATH464.swl.thr3_state;
thread_status[1860] = `IFUPATH465.swl.thr0_state;
thread_status[1861] = `IFUPATH465.swl.thr1_state;
thread_status[1862] = `IFUPATH465.swl.thr2_state;
thread_status[1863] = `IFUPATH465.swl.thr3_state;
thread_status[1864] = `IFUPATH466.swl.thr0_state;
thread_status[1865] = `IFUPATH466.swl.thr1_state;
thread_status[1866] = `IFUPATH466.swl.thr2_state;
thread_status[1867] = `IFUPATH466.swl.thr3_state;
thread_status[1868] = `IFUPATH467.swl.thr0_state;
thread_status[1869] = `IFUPATH467.swl.thr1_state;
thread_status[1870] = `IFUPATH467.swl.thr2_state;
thread_status[1871] = `IFUPATH467.swl.thr3_state;
thread_status[1872] = `IFUPATH468.swl.thr0_state;
thread_status[1873] = `IFUPATH468.swl.thr1_state;
thread_status[1874] = `IFUPATH468.swl.thr2_state;
thread_status[1875] = `IFUPATH468.swl.thr3_state;
thread_status[1876] = `IFUPATH469.swl.thr0_state;
thread_status[1877] = `IFUPATH469.swl.thr1_state;
thread_status[1878] = `IFUPATH469.swl.thr2_state;
thread_status[1879] = `IFUPATH469.swl.thr3_state;
thread_status[1880] = `IFUPATH470.swl.thr0_state;
thread_status[1881] = `IFUPATH470.swl.thr1_state;
thread_status[1882] = `IFUPATH470.swl.thr2_state;
thread_status[1883] = `IFUPATH470.swl.thr3_state;
thread_status[1884] = `IFUPATH471.swl.thr0_state;
thread_status[1885] = `IFUPATH471.swl.thr1_state;
thread_status[1886] = `IFUPATH471.swl.thr2_state;
thread_status[1887] = `IFUPATH471.swl.thr3_state;
thread_status[1888] = `IFUPATH472.swl.thr0_state;
thread_status[1889] = `IFUPATH472.swl.thr1_state;
thread_status[1890] = `IFUPATH472.swl.thr2_state;
thread_status[1891] = `IFUPATH472.swl.thr3_state;
thread_status[1892] = `IFUPATH473.swl.thr0_state;
thread_status[1893] = `IFUPATH473.swl.thr1_state;
thread_status[1894] = `IFUPATH473.swl.thr2_state;
thread_status[1895] = `IFUPATH473.swl.thr3_state;
thread_status[1896] = `IFUPATH474.swl.thr0_state;
thread_status[1897] = `IFUPATH474.swl.thr1_state;
thread_status[1898] = `IFUPATH474.swl.thr2_state;
thread_status[1899] = `IFUPATH474.swl.thr3_state;
thread_status[1900] = `IFUPATH475.swl.thr0_state;
thread_status[1901] = `IFUPATH475.swl.thr1_state;
thread_status[1902] = `IFUPATH475.swl.thr2_state;
thread_status[1903] = `IFUPATH475.swl.thr3_state;
thread_status[1904] = `IFUPATH476.swl.thr0_state;
thread_status[1905] = `IFUPATH476.swl.thr1_state;
thread_status[1906] = `IFUPATH476.swl.thr2_state;
thread_status[1907] = `IFUPATH476.swl.thr3_state;
thread_status[1908] = `IFUPATH477.swl.thr0_state;
thread_status[1909] = `IFUPATH477.swl.thr1_state;
thread_status[1910] = `IFUPATH477.swl.thr2_state;
thread_status[1911] = `IFUPATH477.swl.thr3_state;
thread_status[1912] = `IFUPATH478.swl.thr0_state;
thread_status[1913] = `IFUPATH478.swl.thr1_state;
thread_status[1914] = `IFUPATH478.swl.thr2_state;
thread_status[1915] = `IFUPATH478.swl.thr3_state;
thread_status[1916] = `IFUPATH479.swl.thr0_state;
thread_status[1917] = `IFUPATH479.swl.thr1_state;
thread_status[1918] = `IFUPATH479.swl.thr2_state;
thread_status[1919] = `IFUPATH479.swl.thr3_state;
thread_status[1920] = `IFUPATH480.swl.thr0_state;
thread_status[1921] = `IFUPATH480.swl.thr1_state;
thread_status[1922] = `IFUPATH480.swl.thr2_state;
thread_status[1923] = `IFUPATH480.swl.thr3_state;
thread_status[1924] = `IFUPATH481.swl.thr0_state;
thread_status[1925] = `IFUPATH481.swl.thr1_state;
thread_status[1926] = `IFUPATH481.swl.thr2_state;
thread_status[1927] = `IFUPATH481.swl.thr3_state;
thread_status[1928] = `IFUPATH482.swl.thr0_state;
thread_status[1929] = `IFUPATH482.swl.thr1_state;
thread_status[1930] = `IFUPATH482.swl.thr2_state;
thread_status[1931] = `IFUPATH482.swl.thr3_state;
thread_status[1932] = `IFUPATH483.swl.thr0_state;
thread_status[1933] = `IFUPATH483.swl.thr1_state;
thread_status[1934] = `IFUPATH483.swl.thr2_state;
thread_status[1935] = `IFUPATH483.swl.thr3_state;
thread_status[1936] = `IFUPATH484.swl.thr0_state;
thread_status[1937] = `IFUPATH484.swl.thr1_state;
thread_status[1938] = `IFUPATH484.swl.thr2_state;
thread_status[1939] = `IFUPATH484.swl.thr3_state;
thread_status[1940] = `IFUPATH485.swl.thr0_state;
thread_status[1941] = `IFUPATH485.swl.thr1_state;
thread_status[1942] = `IFUPATH485.swl.thr2_state;
thread_status[1943] = `IFUPATH485.swl.thr3_state;
thread_status[1944] = `IFUPATH486.swl.thr0_state;
thread_status[1945] = `IFUPATH486.swl.thr1_state;
thread_status[1946] = `IFUPATH486.swl.thr2_state;
thread_status[1947] = `IFUPATH486.swl.thr3_state;
thread_status[1948] = `IFUPATH487.swl.thr0_state;
thread_status[1949] = `IFUPATH487.swl.thr1_state;
thread_status[1950] = `IFUPATH487.swl.thr2_state;
thread_status[1951] = `IFUPATH487.swl.thr3_state;
thread_status[1952] = `IFUPATH488.swl.thr0_state;
thread_status[1953] = `IFUPATH488.swl.thr1_state;
thread_status[1954] = `IFUPATH488.swl.thr2_state;
thread_status[1955] = `IFUPATH488.swl.thr3_state;
thread_status[1956] = `IFUPATH489.swl.thr0_state;
thread_status[1957] = `IFUPATH489.swl.thr1_state;
thread_status[1958] = `IFUPATH489.swl.thr2_state;
thread_status[1959] = `IFUPATH489.swl.thr3_state;
thread_status[1960] = `IFUPATH490.swl.thr0_state;
thread_status[1961] = `IFUPATH490.swl.thr1_state;
thread_status[1962] = `IFUPATH490.swl.thr2_state;
thread_status[1963] = `IFUPATH490.swl.thr3_state;
thread_status[1964] = `IFUPATH491.swl.thr0_state;
thread_status[1965] = `IFUPATH491.swl.thr1_state;
thread_status[1966] = `IFUPATH491.swl.thr2_state;
thread_status[1967] = `IFUPATH491.swl.thr3_state;
thread_status[1968] = `IFUPATH492.swl.thr0_state;
thread_status[1969] = `IFUPATH492.swl.thr1_state;
thread_status[1970] = `IFUPATH492.swl.thr2_state;
thread_status[1971] = `IFUPATH492.swl.thr3_state;
thread_status[1972] = `IFUPATH493.swl.thr0_state;
thread_status[1973] = `IFUPATH493.swl.thr1_state;
thread_status[1974] = `IFUPATH493.swl.thr2_state;
thread_status[1975] = `IFUPATH493.swl.thr3_state;
thread_status[1976] = `IFUPATH494.swl.thr0_state;
thread_status[1977] = `IFUPATH494.swl.thr1_state;
thread_status[1978] = `IFUPATH494.swl.thr2_state;
thread_status[1979] = `IFUPATH494.swl.thr3_state;
thread_status[1980] = `IFUPATH495.swl.thr0_state;
thread_status[1981] = `IFUPATH495.swl.thr1_state;
thread_status[1982] = `IFUPATH495.swl.thr2_state;
thread_status[1983] = `IFUPATH495.swl.thr3_state;
thread_status[1984] = `IFUPATH496.swl.thr0_state;
thread_status[1985] = `IFUPATH496.swl.thr1_state;
thread_status[1986] = `IFUPATH496.swl.thr2_state;
thread_status[1987] = `IFUPATH496.swl.thr3_state;
thread_status[1988] = `IFUPATH497.swl.thr0_state;
thread_status[1989] = `IFUPATH497.swl.thr1_state;
thread_status[1990] = `IFUPATH497.swl.thr2_state;
thread_status[1991] = `IFUPATH497.swl.thr3_state;
thread_status[1992] = `IFUPATH498.swl.thr0_state;
thread_status[1993] = `IFUPATH498.swl.thr1_state;
thread_status[1994] = `IFUPATH498.swl.thr2_state;
thread_status[1995] = `IFUPATH498.swl.thr3_state;
thread_status[1996] = `IFUPATH499.swl.thr0_state;
thread_status[1997] = `IFUPATH499.swl.thr1_state;
thread_status[1998] = `IFUPATH499.swl.thr2_state;
thread_status[1999] = `IFUPATH499.swl.thr3_state;
thread_status[2000] = `IFUPATH500.swl.thr0_state;
thread_status[2001] = `IFUPATH500.swl.thr1_state;
thread_status[2002] = `IFUPATH500.swl.thr2_state;
thread_status[2003] = `IFUPATH500.swl.thr3_state;
thread_status[2004] = `IFUPATH501.swl.thr0_state;
thread_status[2005] = `IFUPATH501.swl.thr1_state;
thread_status[2006] = `IFUPATH501.swl.thr2_state;
thread_status[2007] = `IFUPATH501.swl.thr3_state;
thread_status[2008] = `IFUPATH502.swl.thr0_state;
thread_status[2009] = `IFUPATH502.swl.thr1_state;
thread_status[2010] = `IFUPATH502.swl.thr2_state;
thread_status[2011] = `IFUPATH502.swl.thr3_state;
thread_status[2012] = `IFUPATH503.swl.thr0_state;
thread_status[2013] = `IFUPATH503.swl.thr1_state;
thread_status[2014] = `IFUPATH503.swl.thr2_state;
thread_status[2015] = `IFUPATH503.swl.thr3_state;
thread_status[2016] = `IFUPATH504.swl.thr0_state;
thread_status[2017] = `IFUPATH504.swl.thr1_state;
thread_status[2018] = `IFUPATH504.swl.thr2_state;
thread_status[2019] = `IFUPATH504.swl.thr3_state;
thread_status[2020] = `IFUPATH505.swl.thr0_state;
thread_status[2021] = `IFUPATH505.swl.thr1_state;
thread_status[2022] = `IFUPATH505.swl.thr2_state;
thread_status[2023] = `IFUPATH505.swl.thr3_state;
thread_status[2024] = `IFUPATH506.swl.thr0_state;
thread_status[2025] = `IFUPATH506.swl.thr1_state;
thread_status[2026] = `IFUPATH506.swl.thr2_state;
thread_status[2027] = `IFUPATH506.swl.thr3_state;
thread_status[2028] = `IFUPATH507.swl.thr0_state;
thread_status[2029] = `IFUPATH507.swl.thr1_state;
thread_status[2030] = `IFUPATH507.swl.thr2_state;
thread_status[2031] = `IFUPATH507.swl.thr3_state;
thread_status[2032] = `IFUPATH508.swl.thr0_state;
thread_status[2033] = `IFUPATH508.swl.thr1_state;
thread_status[2034] = `IFUPATH508.swl.thr2_state;
thread_status[2035] = `IFUPATH508.swl.thr3_state;
thread_status[2036] = `IFUPATH509.swl.thr0_state;
thread_status[2037] = `IFUPATH509.swl.thr1_state;
thread_status[2038] = `IFUPATH509.swl.thr2_state;
thread_status[2039] = `IFUPATH509.swl.thr3_state;
thread_status[2040] = `IFUPATH510.swl.thr0_state;
thread_status[2041] = `IFUPATH510.swl.thr1_state;
thread_status[2042] = `IFUPATH510.swl.thr2_state;
thread_status[2043] = `IFUPATH510.swl.thr3_state;
thread_status[2044] = `IFUPATH511.swl.thr0_state;
thread_status[2045] = `IFUPATH511.swl.thr1_state;
thread_status[2046] = `IFUPATH511.swl.thr2_state;
thread_status[2047] = `IFUPATH511.swl.thr3_state;
thread_status[2048] = `IFUPATH512.swl.thr0_state;
thread_status[2049] = `IFUPATH512.swl.thr1_state;
thread_status[2050] = `IFUPATH512.swl.thr2_state;
thread_status[2051] = `IFUPATH512.swl.thr3_state;
thread_status[2052] = `IFUPATH513.swl.thr0_state;
thread_status[2053] = `IFUPATH513.swl.thr1_state;
thread_status[2054] = `IFUPATH513.swl.thr2_state;
thread_status[2055] = `IFUPATH513.swl.thr3_state;
thread_status[2056] = `IFUPATH514.swl.thr0_state;
thread_status[2057] = `IFUPATH514.swl.thr1_state;
thread_status[2058] = `IFUPATH514.swl.thr2_state;
thread_status[2059] = `IFUPATH514.swl.thr3_state;
thread_status[2060] = `IFUPATH515.swl.thr0_state;
thread_status[2061] = `IFUPATH515.swl.thr1_state;
thread_status[2062] = `IFUPATH515.swl.thr2_state;
thread_status[2063] = `IFUPATH515.swl.thr3_state;
thread_status[2064] = `IFUPATH516.swl.thr0_state;
thread_status[2065] = `IFUPATH516.swl.thr1_state;
thread_status[2066] = `IFUPATH516.swl.thr2_state;
thread_status[2067] = `IFUPATH516.swl.thr3_state;
thread_status[2068] = `IFUPATH517.swl.thr0_state;
thread_status[2069] = `IFUPATH517.swl.thr1_state;
thread_status[2070] = `IFUPATH517.swl.thr2_state;
thread_status[2071] = `IFUPATH517.swl.thr3_state;
thread_status[2072] = `IFUPATH518.swl.thr0_state;
thread_status[2073] = `IFUPATH518.swl.thr1_state;
thread_status[2074] = `IFUPATH518.swl.thr2_state;
thread_status[2075] = `IFUPATH518.swl.thr3_state;
thread_status[2076] = `IFUPATH519.swl.thr0_state;
thread_status[2077] = `IFUPATH519.swl.thr1_state;
thread_status[2078] = `IFUPATH519.swl.thr2_state;
thread_status[2079] = `IFUPATH519.swl.thr3_state;
thread_status[2080] = `IFUPATH520.swl.thr0_state;
thread_status[2081] = `IFUPATH520.swl.thr1_state;
thread_status[2082] = `IFUPATH520.swl.thr2_state;
thread_status[2083] = `IFUPATH520.swl.thr3_state;
thread_status[2084] = `IFUPATH521.swl.thr0_state;
thread_status[2085] = `IFUPATH521.swl.thr1_state;
thread_status[2086] = `IFUPATH521.swl.thr2_state;
thread_status[2087] = `IFUPATH521.swl.thr3_state;
thread_status[2088] = `IFUPATH522.swl.thr0_state;
thread_status[2089] = `IFUPATH522.swl.thr1_state;
thread_status[2090] = `IFUPATH522.swl.thr2_state;
thread_status[2091] = `IFUPATH522.swl.thr3_state;
thread_status[2092] = `IFUPATH523.swl.thr0_state;
thread_status[2093] = `IFUPATH523.swl.thr1_state;
thread_status[2094] = `IFUPATH523.swl.thr2_state;
thread_status[2095] = `IFUPATH523.swl.thr3_state;
thread_status[2096] = `IFUPATH524.swl.thr0_state;
thread_status[2097] = `IFUPATH524.swl.thr1_state;
thread_status[2098] = `IFUPATH524.swl.thr2_state;
thread_status[2099] = `IFUPATH524.swl.thr3_state;
thread_status[2100] = `IFUPATH525.swl.thr0_state;
thread_status[2101] = `IFUPATH525.swl.thr1_state;
thread_status[2102] = `IFUPATH525.swl.thr2_state;
thread_status[2103] = `IFUPATH525.swl.thr3_state;
thread_status[2104] = `IFUPATH526.swl.thr0_state;
thread_status[2105] = `IFUPATH526.swl.thr1_state;
thread_status[2106] = `IFUPATH526.swl.thr2_state;
thread_status[2107] = `IFUPATH526.swl.thr3_state;
thread_status[2108] = `IFUPATH527.swl.thr0_state;
thread_status[2109] = `IFUPATH527.swl.thr1_state;
thread_status[2110] = `IFUPATH527.swl.thr2_state;
thread_status[2111] = `IFUPATH527.swl.thr3_state;
thread_status[2112] = `IFUPATH528.swl.thr0_state;
thread_status[2113] = `IFUPATH528.swl.thr1_state;
thread_status[2114] = `IFUPATH528.swl.thr2_state;
thread_status[2115] = `IFUPATH528.swl.thr3_state;
thread_status[2116] = `IFUPATH529.swl.thr0_state;
thread_status[2117] = `IFUPATH529.swl.thr1_state;
thread_status[2118] = `IFUPATH529.swl.thr2_state;
thread_status[2119] = `IFUPATH529.swl.thr3_state;
thread_status[2120] = `IFUPATH530.swl.thr0_state;
thread_status[2121] = `IFUPATH530.swl.thr1_state;
thread_status[2122] = `IFUPATH530.swl.thr2_state;
thread_status[2123] = `IFUPATH530.swl.thr3_state;
thread_status[2124] = `IFUPATH531.swl.thr0_state;
thread_status[2125] = `IFUPATH531.swl.thr1_state;
thread_status[2126] = `IFUPATH531.swl.thr2_state;
thread_status[2127] = `IFUPATH531.swl.thr3_state;
thread_status[2128] = `IFUPATH532.swl.thr0_state;
thread_status[2129] = `IFUPATH532.swl.thr1_state;
thread_status[2130] = `IFUPATH532.swl.thr2_state;
thread_status[2131] = `IFUPATH532.swl.thr3_state;
thread_status[2132] = `IFUPATH533.swl.thr0_state;
thread_status[2133] = `IFUPATH533.swl.thr1_state;
thread_status[2134] = `IFUPATH533.swl.thr2_state;
thread_status[2135] = `IFUPATH533.swl.thr3_state;
thread_status[2136] = `IFUPATH534.swl.thr0_state;
thread_status[2137] = `IFUPATH534.swl.thr1_state;
thread_status[2138] = `IFUPATH534.swl.thr2_state;
thread_status[2139] = `IFUPATH534.swl.thr3_state;
thread_status[2140] = `IFUPATH535.swl.thr0_state;
thread_status[2141] = `IFUPATH535.swl.thr1_state;
thread_status[2142] = `IFUPATH535.swl.thr2_state;
thread_status[2143] = `IFUPATH535.swl.thr3_state;
thread_status[2144] = `IFUPATH536.swl.thr0_state;
thread_status[2145] = `IFUPATH536.swl.thr1_state;
thread_status[2146] = `IFUPATH536.swl.thr2_state;
thread_status[2147] = `IFUPATH536.swl.thr3_state;
thread_status[2148] = `IFUPATH537.swl.thr0_state;
thread_status[2149] = `IFUPATH537.swl.thr1_state;
thread_status[2150] = `IFUPATH537.swl.thr2_state;
thread_status[2151] = `IFUPATH537.swl.thr3_state;
thread_status[2152] = `IFUPATH538.swl.thr0_state;
thread_status[2153] = `IFUPATH538.swl.thr1_state;
thread_status[2154] = `IFUPATH538.swl.thr2_state;
thread_status[2155] = `IFUPATH538.swl.thr3_state;
thread_status[2156] = `IFUPATH539.swl.thr0_state;
thread_status[2157] = `IFUPATH539.swl.thr1_state;
thread_status[2158] = `IFUPATH539.swl.thr2_state;
thread_status[2159] = `IFUPATH539.swl.thr3_state;
thread_status[2160] = `IFUPATH540.swl.thr0_state;
thread_status[2161] = `IFUPATH540.swl.thr1_state;
thread_status[2162] = `IFUPATH540.swl.thr2_state;
thread_status[2163] = `IFUPATH540.swl.thr3_state;
thread_status[2164] = `IFUPATH541.swl.thr0_state;
thread_status[2165] = `IFUPATH541.swl.thr1_state;
thread_status[2166] = `IFUPATH541.swl.thr2_state;
thread_status[2167] = `IFUPATH541.swl.thr3_state;
thread_status[2168] = `IFUPATH542.swl.thr0_state;
thread_status[2169] = `IFUPATH542.swl.thr1_state;
thread_status[2170] = `IFUPATH542.swl.thr2_state;
thread_status[2171] = `IFUPATH542.swl.thr3_state;
thread_status[2172] = `IFUPATH543.swl.thr0_state;
thread_status[2173] = `IFUPATH543.swl.thr1_state;
thread_status[2174] = `IFUPATH543.swl.thr2_state;
thread_status[2175] = `IFUPATH543.swl.thr3_state;
thread_status[2176] = `IFUPATH544.swl.thr0_state;
thread_status[2177] = `IFUPATH544.swl.thr1_state;
thread_status[2178] = `IFUPATH544.swl.thr2_state;
thread_status[2179] = `IFUPATH544.swl.thr3_state;
thread_status[2180] = `IFUPATH545.swl.thr0_state;
thread_status[2181] = `IFUPATH545.swl.thr1_state;
thread_status[2182] = `IFUPATH545.swl.thr2_state;
thread_status[2183] = `IFUPATH545.swl.thr3_state;
thread_status[2184] = `IFUPATH546.swl.thr0_state;
thread_status[2185] = `IFUPATH546.swl.thr1_state;
thread_status[2186] = `IFUPATH546.swl.thr2_state;
thread_status[2187] = `IFUPATH546.swl.thr3_state;
thread_status[2188] = `IFUPATH547.swl.thr0_state;
thread_status[2189] = `IFUPATH547.swl.thr1_state;
thread_status[2190] = `IFUPATH547.swl.thr2_state;
thread_status[2191] = `IFUPATH547.swl.thr3_state;
thread_status[2192] = `IFUPATH548.swl.thr0_state;
thread_status[2193] = `IFUPATH548.swl.thr1_state;
thread_status[2194] = `IFUPATH548.swl.thr2_state;
thread_status[2195] = `IFUPATH548.swl.thr3_state;
thread_status[2196] = `IFUPATH549.swl.thr0_state;
thread_status[2197] = `IFUPATH549.swl.thr1_state;
thread_status[2198] = `IFUPATH549.swl.thr2_state;
thread_status[2199] = `IFUPATH549.swl.thr3_state;
thread_status[2200] = `IFUPATH550.swl.thr0_state;
thread_status[2201] = `IFUPATH550.swl.thr1_state;
thread_status[2202] = `IFUPATH550.swl.thr2_state;
thread_status[2203] = `IFUPATH550.swl.thr3_state;
thread_status[2204] = `IFUPATH551.swl.thr0_state;
thread_status[2205] = `IFUPATH551.swl.thr1_state;
thread_status[2206] = `IFUPATH551.swl.thr2_state;
thread_status[2207] = `IFUPATH551.swl.thr3_state;
thread_status[2208] = `IFUPATH552.swl.thr0_state;
thread_status[2209] = `IFUPATH552.swl.thr1_state;
thread_status[2210] = `IFUPATH552.swl.thr2_state;
thread_status[2211] = `IFUPATH552.swl.thr3_state;
thread_status[2212] = `IFUPATH553.swl.thr0_state;
thread_status[2213] = `IFUPATH553.swl.thr1_state;
thread_status[2214] = `IFUPATH553.swl.thr2_state;
thread_status[2215] = `IFUPATH553.swl.thr3_state;
thread_status[2216] = `IFUPATH554.swl.thr0_state;
thread_status[2217] = `IFUPATH554.swl.thr1_state;
thread_status[2218] = `IFUPATH554.swl.thr2_state;
thread_status[2219] = `IFUPATH554.swl.thr3_state;
thread_status[2220] = `IFUPATH555.swl.thr0_state;
thread_status[2221] = `IFUPATH555.swl.thr1_state;
thread_status[2222] = `IFUPATH555.swl.thr2_state;
thread_status[2223] = `IFUPATH555.swl.thr3_state;
thread_status[2224] = `IFUPATH556.swl.thr0_state;
thread_status[2225] = `IFUPATH556.swl.thr1_state;
thread_status[2226] = `IFUPATH556.swl.thr2_state;
thread_status[2227] = `IFUPATH556.swl.thr3_state;
thread_status[2228] = `IFUPATH557.swl.thr0_state;
thread_status[2229] = `IFUPATH557.swl.thr1_state;
thread_status[2230] = `IFUPATH557.swl.thr2_state;
thread_status[2231] = `IFUPATH557.swl.thr3_state;
thread_status[2232] = `IFUPATH558.swl.thr0_state;
thread_status[2233] = `IFUPATH558.swl.thr1_state;
thread_status[2234] = `IFUPATH558.swl.thr2_state;
thread_status[2235] = `IFUPATH558.swl.thr3_state;
thread_status[2236] = `IFUPATH559.swl.thr0_state;
thread_status[2237] = `IFUPATH559.swl.thr1_state;
thread_status[2238] = `IFUPATH559.swl.thr2_state;
thread_status[2239] = `IFUPATH559.swl.thr3_state;
thread_status[2240] = `IFUPATH560.swl.thr0_state;
thread_status[2241] = `IFUPATH560.swl.thr1_state;
thread_status[2242] = `IFUPATH560.swl.thr2_state;
thread_status[2243] = `IFUPATH560.swl.thr3_state;
thread_status[2244] = `IFUPATH561.swl.thr0_state;
thread_status[2245] = `IFUPATH561.swl.thr1_state;
thread_status[2246] = `IFUPATH561.swl.thr2_state;
thread_status[2247] = `IFUPATH561.swl.thr3_state;
thread_status[2248] = `IFUPATH562.swl.thr0_state;
thread_status[2249] = `IFUPATH562.swl.thr1_state;
thread_status[2250] = `IFUPATH562.swl.thr2_state;
thread_status[2251] = `IFUPATH562.swl.thr3_state;
thread_status[2252] = `IFUPATH563.swl.thr0_state;
thread_status[2253] = `IFUPATH563.swl.thr1_state;
thread_status[2254] = `IFUPATH563.swl.thr2_state;
thread_status[2255] = `IFUPATH563.swl.thr3_state;
thread_status[2256] = `IFUPATH564.swl.thr0_state;
thread_status[2257] = `IFUPATH564.swl.thr1_state;
thread_status[2258] = `IFUPATH564.swl.thr2_state;
thread_status[2259] = `IFUPATH564.swl.thr3_state;
thread_status[2260] = `IFUPATH565.swl.thr0_state;
thread_status[2261] = `IFUPATH565.swl.thr1_state;
thread_status[2262] = `IFUPATH565.swl.thr2_state;
thread_status[2263] = `IFUPATH565.swl.thr3_state;
thread_status[2264] = `IFUPATH566.swl.thr0_state;
thread_status[2265] = `IFUPATH566.swl.thr1_state;
thread_status[2266] = `IFUPATH566.swl.thr2_state;
thread_status[2267] = `IFUPATH566.swl.thr3_state;
thread_status[2268] = `IFUPATH567.swl.thr0_state;
thread_status[2269] = `IFUPATH567.swl.thr1_state;
thread_status[2270] = `IFUPATH567.swl.thr2_state;
thread_status[2271] = `IFUPATH567.swl.thr3_state;
thread_status[2272] = `IFUPATH568.swl.thr0_state;
thread_status[2273] = `IFUPATH568.swl.thr1_state;
thread_status[2274] = `IFUPATH568.swl.thr2_state;
thread_status[2275] = `IFUPATH568.swl.thr3_state;
thread_status[2276] = `IFUPATH569.swl.thr0_state;
thread_status[2277] = `IFUPATH569.swl.thr1_state;
thread_status[2278] = `IFUPATH569.swl.thr2_state;
thread_status[2279] = `IFUPATH569.swl.thr3_state;
thread_status[2280] = `IFUPATH570.swl.thr0_state;
thread_status[2281] = `IFUPATH570.swl.thr1_state;
thread_status[2282] = `IFUPATH570.swl.thr2_state;
thread_status[2283] = `IFUPATH570.swl.thr3_state;
thread_status[2284] = `IFUPATH571.swl.thr0_state;
thread_status[2285] = `IFUPATH571.swl.thr1_state;
thread_status[2286] = `IFUPATH571.swl.thr2_state;
thread_status[2287] = `IFUPATH571.swl.thr3_state;
thread_status[2288] = `IFUPATH572.swl.thr0_state;
thread_status[2289] = `IFUPATH572.swl.thr1_state;
thread_status[2290] = `IFUPATH572.swl.thr2_state;
thread_status[2291] = `IFUPATH572.swl.thr3_state;
thread_status[2292] = `IFUPATH573.swl.thr0_state;
thread_status[2293] = `IFUPATH573.swl.thr1_state;
thread_status[2294] = `IFUPATH573.swl.thr2_state;
thread_status[2295] = `IFUPATH573.swl.thr3_state;
thread_status[2296] = `IFUPATH574.swl.thr0_state;
thread_status[2297] = `IFUPATH574.swl.thr1_state;
thread_status[2298] = `IFUPATH574.swl.thr2_state;
thread_status[2299] = `IFUPATH574.swl.thr3_state;
thread_status[2300] = `IFUPATH575.swl.thr0_state;
thread_status[2301] = `IFUPATH575.swl.thr1_state;
thread_status[2302] = `IFUPATH575.swl.thr2_state;
thread_status[2303] = `IFUPATH575.swl.thr3_state;
thread_status[2304] = `IFUPATH576.swl.thr0_state;
thread_status[2305] = `IFUPATH576.swl.thr1_state;
thread_status[2306] = `IFUPATH576.swl.thr2_state;
thread_status[2307] = `IFUPATH576.swl.thr3_state;
thread_status[2308] = `IFUPATH577.swl.thr0_state;
thread_status[2309] = `IFUPATH577.swl.thr1_state;
thread_status[2310] = `IFUPATH577.swl.thr2_state;
thread_status[2311] = `IFUPATH577.swl.thr3_state;
thread_status[2312] = `IFUPATH578.swl.thr0_state;
thread_status[2313] = `IFUPATH578.swl.thr1_state;
thread_status[2314] = `IFUPATH578.swl.thr2_state;
thread_status[2315] = `IFUPATH578.swl.thr3_state;
thread_status[2316] = `IFUPATH579.swl.thr0_state;
thread_status[2317] = `IFUPATH579.swl.thr1_state;
thread_status[2318] = `IFUPATH579.swl.thr2_state;
thread_status[2319] = `IFUPATH579.swl.thr3_state;
thread_status[2320] = `IFUPATH580.swl.thr0_state;
thread_status[2321] = `IFUPATH580.swl.thr1_state;
thread_status[2322] = `IFUPATH580.swl.thr2_state;
thread_status[2323] = `IFUPATH580.swl.thr3_state;
thread_status[2324] = `IFUPATH581.swl.thr0_state;
thread_status[2325] = `IFUPATH581.swl.thr1_state;
thread_status[2326] = `IFUPATH581.swl.thr2_state;
thread_status[2327] = `IFUPATH581.swl.thr3_state;
thread_status[2328] = `IFUPATH582.swl.thr0_state;
thread_status[2329] = `IFUPATH582.swl.thr1_state;
thread_status[2330] = `IFUPATH582.swl.thr2_state;
thread_status[2331] = `IFUPATH582.swl.thr3_state;
thread_status[2332] = `IFUPATH583.swl.thr0_state;
thread_status[2333] = `IFUPATH583.swl.thr1_state;
thread_status[2334] = `IFUPATH583.swl.thr2_state;
thread_status[2335] = `IFUPATH583.swl.thr3_state;
thread_status[2336] = `IFUPATH584.swl.thr0_state;
thread_status[2337] = `IFUPATH584.swl.thr1_state;
thread_status[2338] = `IFUPATH584.swl.thr2_state;
thread_status[2339] = `IFUPATH584.swl.thr3_state;
thread_status[2340] = `IFUPATH585.swl.thr0_state;
thread_status[2341] = `IFUPATH585.swl.thr1_state;
thread_status[2342] = `IFUPATH585.swl.thr2_state;
thread_status[2343] = `IFUPATH585.swl.thr3_state;
thread_status[2344] = `IFUPATH586.swl.thr0_state;
thread_status[2345] = `IFUPATH586.swl.thr1_state;
thread_status[2346] = `IFUPATH586.swl.thr2_state;
thread_status[2347] = `IFUPATH586.swl.thr3_state;
thread_status[2348] = `IFUPATH587.swl.thr0_state;
thread_status[2349] = `IFUPATH587.swl.thr1_state;
thread_status[2350] = `IFUPATH587.swl.thr2_state;
thread_status[2351] = `IFUPATH587.swl.thr3_state;
thread_status[2352] = `IFUPATH588.swl.thr0_state;
thread_status[2353] = `IFUPATH588.swl.thr1_state;
thread_status[2354] = `IFUPATH588.swl.thr2_state;
thread_status[2355] = `IFUPATH588.swl.thr3_state;
thread_status[2356] = `IFUPATH589.swl.thr0_state;
thread_status[2357] = `IFUPATH589.swl.thr1_state;
thread_status[2358] = `IFUPATH589.swl.thr2_state;
thread_status[2359] = `IFUPATH589.swl.thr3_state;
thread_status[2360] = `IFUPATH590.swl.thr0_state;
thread_status[2361] = `IFUPATH590.swl.thr1_state;
thread_status[2362] = `IFUPATH590.swl.thr2_state;
thread_status[2363] = `IFUPATH590.swl.thr3_state;
thread_status[2364] = `IFUPATH591.swl.thr0_state;
thread_status[2365] = `IFUPATH591.swl.thr1_state;
thread_status[2366] = `IFUPATH591.swl.thr2_state;
thread_status[2367] = `IFUPATH591.swl.thr3_state;
thread_status[2368] = `IFUPATH592.swl.thr0_state;
thread_status[2369] = `IFUPATH592.swl.thr1_state;
thread_status[2370] = `IFUPATH592.swl.thr2_state;
thread_status[2371] = `IFUPATH592.swl.thr3_state;
thread_status[2372] = `IFUPATH593.swl.thr0_state;
thread_status[2373] = `IFUPATH593.swl.thr1_state;
thread_status[2374] = `IFUPATH593.swl.thr2_state;
thread_status[2375] = `IFUPATH593.swl.thr3_state;
thread_status[2376] = `IFUPATH594.swl.thr0_state;
thread_status[2377] = `IFUPATH594.swl.thr1_state;
thread_status[2378] = `IFUPATH594.swl.thr2_state;
thread_status[2379] = `IFUPATH594.swl.thr3_state;
thread_status[2380] = `IFUPATH595.swl.thr0_state;
thread_status[2381] = `IFUPATH595.swl.thr1_state;
thread_status[2382] = `IFUPATH595.swl.thr2_state;
thread_status[2383] = `IFUPATH595.swl.thr3_state;
thread_status[2384] = `IFUPATH596.swl.thr0_state;
thread_status[2385] = `IFUPATH596.swl.thr1_state;
thread_status[2386] = `IFUPATH596.swl.thr2_state;
thread_status[2387] = `IFUPATH596.swl.thr3_state;
thread_status[2388] = `IFUPATH597.swl.thr0_state;
thread_status[2389] = `IFUPATH597.swl.thr1_state;
thread_status[2390] = `IFUPATH597.swl.thr2_state;
thread_status[2391] = `IFUPATH597.swl.thr3_state;
thread_status[2392] = `IFUPATH598.swl.thr0_state;
thread_status[2393] = `IFUPATH598.swl.thr1_state;
thread_status[2394] = `IFUPATH598.swl.thr2_state;
thread_status[2395] = `IFUPATH598.swl.thr3_state;
thread_status[2396] = `IFUPATH599.swl.thr0_state;
thread_status[2397] = `IFUPATH599.swl.thr1_state;
thread_status[2398] = `IFUPATH599.swl.thr2_state;
thread_status[2399] = `IFUPATH599.swl.thr3_state;
thread_status[2400] = `IFUPATH600.swl.thr0_state;
thread_status[2401] = `IFUPATH600.swl.thr1_state;
thread_status[2402] = `IFUPATH600.swl.thr2_state;
thread_status[2403] = `IFUPATH600.swl.thr3_state;
thread_status[2404] = `IFUPATH601.swl.thr0_state;
thread_status[2405] = `IFUPATH601.swl.thr1_state;
thread_status[2406] = `IFUPATH601.swl.thr2_state;
thread_status[2407] = `IFUPATH601.swl.thr3_state;
thread_status[2408] = `IFUPATH602.swl.thr0_state;
thread_status[2409] = `IFUPATH602.swl.thr1_state;
thread_status[2410] = `IFUPATH602.swl.thr2_state;
thread_status[2411] = `IFUPATH602.swl.thr3_state;
thread_status[2412] = `IFUPATH603.swl.thr0_state;
thread_status[2413] = `IFUPATH603.swl.thr1_state;
thread_status[2414] = `IFUPATH603.swl.thr2_state;
thread_status[2415] = `IFUPATH603.swl.thr3_state;
thread_status[2416] = `IFUPATH604.swl.thr0_state;
thread_status[2417] = `IFUPATH604.swl.thr1_state;
thread_status[2418] = `IFUPATH604.swl.thr2_state;
thread_status[2419] = `IFUPATH604.swl.thr3_state;
thread_status[2420] = `IFUPATH605.swl.thr0_state;
thread_status[2421] = `IFUPATH605.swl.thr1_state;
thread_status[2422] = `IFUPATH605.swl.thr2_state;
thread_status[2423] = `IFUPATH605.swl.thr3_state;
thread_status[2424] = `IFUPATH606.swl.thr0_state;
thread_status[2425] = `IFUPATH606.swl.thr1_state;
thread_status[2426] = `IFUPATH606.swl.thr2_state;
thread_status[2427] = `IFUPATH606.swl.thr3_state;
thread_status[2428] = `IFUPATH607.swl.thr0_state;
thread_status[2429] = `IFUPATH607.swl.thr1_state;
thread_status[2430] = `IFUPATH607.swl.thr2_state;
thread_status[2431] = `IFUPATH607.swl.thr3_state;
thread_status[2432] = `IFUPATH608.swl.thr0_state;
thread_status[2433] = `IFUPATH608.swl.thr1_state;
thread_status[2434] = `IFUPATH608.swl.thr2_state;
thread_status[2435] = `IFUPATH608.swl.thr3_state;
thread_status[2436] = `IFUPATH609.swl.thr0_state;
thread_status[2437] = `IFUPATH609.swl.thr1_state;
thread_status[2438] = `IFUPATH609.swl.thr2_state;
thread_status[2439] = `IFUPATH609.swl.thr3_state;
thread_status[2440] = `IFUPATH610.swl.thr0_state;
thread_status[2441] = `IFUPATH610.swl.thr1_state;
thread_status[2442] = `IFUPATH610.swl.thr2_state;
thread_status[2443] = `IFUPATH610.swl.thr3_state;
thread_status[2444] = `IFUPATH611.swl.thr0_state;
thread_status[2445] = `IFUPATH611.swl.thr1_state;
thread_status[2446] = `IFUPATH611.swl.thr2_state;
thread_status[2447] = `IFUPATH611.swl.thr3_state;
thread_status[2448] = `IFUPATH612.swl.thr0_state;
thread_status[2449] = `IFUPATH612.swl.thr1_state;
thread_status[2450] = `IFUPATH612.swl.thr2_state;
thread_status[2451] = `IFUPATH612.swl.thr3_state;
thread_status[2452] = `IFUPATH613.swl.thr0_state;
thread_status[2453] = `IFUPATH613.swl.thr1_state;
thread_status[2454] = `IFUPATH613.swl.thr2_state;
thread_status[2455] = `IFUPATH613.swl.thr3_state;
thread_status[2456] = `IFUPATH614.swl.thr0_state;
thread_status[2457] = `IFUPATH614.swl.thr1_state;
thread_status[2458] = `IFUPATH614.swl.thr2_state;
thread_status[2459] = `IFUPATH614.swl.thr3_state;
thread_status[2460] = `IFUPATH615.swl.thr0_state;
thread_status[2461] = `IFUPATH615.swl.thr1_state;
thread_status[2462] = `IFUPATH615.swl.thr2_state;
thread_status[2463] = `IFUPATH615.swl.thr3_state;
thread_status[2464] = `IFUPATH616.swl.thr0_state;
thread_status[2465] = `IFUPATH616.swl.thr1_state;
thread_status[2466] = `IFUPATH616.swl.thr2_state;
thread_status[2467] = `IFUPATH616.swl.thr3_state;
thread_status[2468] = `IFUPATH617.swl.thr0_state;
thread_status[2469] = `IFUPATH617.swl.thr1_state;
thread_status[2470] = `IFUPATH617.swl.thr2_state;
thread_status[2471] = `IFUPATH617.swl.thr3_state;
thread_status[2472] = `IFUPATH618.swl.thr0_state;
thread_status[2473] = `IFUPATH618.swl.thr1_state;
thread_status[2474] = `IFUPATH618.swl.thr2_state;
thread_status[2475] = `IFUPATH618.swl.thr3_state;
thread_status[2476] = `IFUPATH619.swl.thr0_state;
thread_status[2477] = `IFUPATH619.swl.thr1_state;
thread_status[2478] = `IFUPATH619.swl.thr2_state;
thread_status[2479] = `IFUPATH619.swl.thr3_state;
thread_status[2480] = `IFUPATH620.swl.thr0_state;
thread_status[2481] = `IFUPATH620.swl.thr1_state;
thread_status[2482] = `IFUPATH620.swl.thr2_state;
thread_status[2483] = `IFUPATH620.swl.thr3_state;
thread_status[2484] = `IFUPATH621.swl.thr0_state;
thread_status[2485] = `IFUPATH621.swl.thr1_state;
thread_status[2486] = `IFUPATH621.swl.thr2_state;
thread_status[2487] = `IFUPATH621.swl.thr3_state;
thread_status[2488] = `IFUPATH622.swl.thr0_state;
thread_status[2489] = `IFUPATH622.swl.thr1_state;
thread_status[2490] = `IFUPATH622.swl.thr2_state;
thread_status[2491] = `IFUPATH622.swl.thr3_state;
thread_status[2492] = `IFUPATH623.swl.thr0_state;
thread_status[2493] = `IFUPATH623.swl.thr1_state;
thread_status[2494] = `IFUPATH623.swl.thr2_state;
thread_status[2495] = `IFUPATH623.swl.thr3_state;
thread_status[2496] = `IFUPATH624.swl.thr0_state;
thread_status[2497] = `IFUPATH624.swl.thr1_state;
thread_status[2498] = `IFUPATH624.swl.thr2_state;
thread_status[2499] = `IFUPATH624.swl.thr3_state;
thread_status[2500] = `IFUPATH625.swl.thr0_state;
thread_status[2501] = `IFUPATH625.swl.thr1_state;
thread_status[2502] = `IFUPATH625.swl.thr2_state;
thread_status[2503] = `IFUPATH625.swl.thr3_state;
thread_status[2504] = `IFUPATH626.swl.thr0_state;
thread_status[2505] = `IFUPATH626.swl.thr1_state;
thread_status[2506] = `IFUPATH626.swl.thr2_state;
thread_status[2507] = `IFUPATH626.swl.thr3_state;
thread_status[2508] = `IFUPATH627.swl.thr0_state;
thread_status[2509] = `IFUPATH627.swl.thr1_state;
thread_status[2510] = `IFUPATH627.swl.thr2_state;
thread_status[2511] = `IFUPATH627.swl.thr3_state;
thread_status[2512] = `IFUPATH628.swl.thr0_state;
thread_status[2513] = `IFUPATH628.swl.thr1_state;
thread_status[2514] = `IFUPATH628.swl.thr2_state;
thread_status[2515] = `IFUPATH628.swl.thr3_state;
thread_status[2516] = `IFUPATH629.swl.thr0_state;
thread_status[2517] = `IFUPATH629.swl.thr1_state;
thread_status[2518] = `IFUPATH629.swl.thr2_state;
thread_status[2519] = `IFUPATH629.swl.thr3_state;
thread_status[2520] = `IFUPATH630.swl.thr0_state;
thread_status[2521] = `IFUPATH630.swl.thr1_state;
thread_status[2522] = `IFUPATH630.swl.thr2_state;
thread_status[2523] = `IFUPATH630.swl.thr3_state;
thread_status[2524] = `IFUPATH631.swl.thr0_state;
thread_status[2525] = `IFUPATH631.swl.thr1_state;
thread_status[2526] = `IFUPATH631.swl.thr2_state;
thread_status[2527] = `IFUPATH631.swl.thr3_state;
thread_status[2528] = `IFUPATH632.swl.thr0_state;
thread_status[2529] = `IFUPATH632.swl.thr1_state;
thread_status[2530] = `IFUPATH632.swl.thr2_state;
thread_status[2531] = `IFUPATH632.swl.thr3_state;
thread_status[2532] = `IFUPATH633.swl.thr0_state;
thread_status[2533] = `IFUPATH633.swl.thr1_state;
thread_status[2534] = `IFUPATH633.swl.thr2_state;
thread_status[2535] = `IFUPATH633.swl.thr3_state;
thread_status[2536] = `IFUPATH634.swl.thr0_state;
thread_status[2537] = `IFUPATH634.swl.thr1_state;
thread_status[2538] = `IFUPATH634.swl.thr2_state;
thread_status[2539] = `IFUPATH634.swl.thr3_state;
thread_status[2540] = `IFUPATH635.swl.thr0_state;
thread_status[2541] = `IFUPATH635.swl.thr1_state;
thread_status[2542] = `IFUPATH635.swl.thr2_state;
thread_status[2543] = `IFUPATH635.swl.thr3_state;
thread_status[2544] = `IFUPATH636.swl.thr0_state;
thread_status[2545] = `IFUPATH636.swl.thr1_state;
thread_status[2546] = `IFUPATH636.swl.thr2_state;
thread_status[2547] = `IFUPATH636.swl.thr3_state;
thread_status[2548] = `IFUPATH637.swl.thr0_state;
thread_status[2549] = `IFUPATH637.swl.thr1_state;
thread_status[2550] = `IFUPATH637.swl.thr2_state;
thread_status[2551] = `IFUPATH637.swl.thr3_state;
thread_status[2552] = `IFUPATH638.swl.thr0_state;
thread_status[2553] = `IFUPATH638.swl.thr1_state;
thread_status[2554] = `IFUPATH638.swl.thr2_state;
thread_status[2555] = `IFUPATH638.swl.thr3_state;
thread_status[2556] = `IFUPATH639.swl.thr0_state;
thread_status[2557] = `IFUPATH639.swl.thr1_state;
thread_status[2558] = `IFUPATH639.swl.thr2_state;
thread_status[2559] = `IFUPATH639.swl.thr3_state;
thread_status[2560] = `IFUPATH640.swl.thr0_state;
thread_status[2561] = `IFUPATH640.swl.thr1_state;
thread_status[2562] = `IFUPATH640.swl.thr2_state;
thread_status[2563] = `IFUPATH640.swl.thr3_state;
thread_status[2564] = `IFUPATH641.swl.thr0_state;
thread_status[2565] = `IFUPATH641.swl.thr1_state;
thread_status[2566] = `IFUPATH641.swl.thr2_state;
thread_status[2567] = `IFUPATH641.swl.thr3_state;
thread_status[2568] = `IFUPATH642.swl.thr0_state;
thread_status[2569] = `IFUPATH642.swl.thr1_state;
thread_status[2570] = `IFUPATH642.swl.thr2_state;
thread_status[2571] = `IFUPATH642.swl.thr3_state;
thread_status[2572] = `IFUPATH643.swl.thr0_state;
thread_status[2573] = `IFUPATH643.swl.thr1_state;
thread_status[2574] = `IFUPATH643.swl.thr2_state;
thread_status[2575] = `IFUPATH643.swl.thr3_state;
thread_status[2576] = `IFUPATH644.swl.thr0_state;
thread_status[2577] = `IFUPATH644.swl.thr1_state;
thread_status[2578] = `IFUPATH644.swl.thr2_state;
thread_status[2579] = `IFUPATH644.swl.thr3_state;
thread_status[2580] = `IFUPATH645.swl.thr0_state;
thread_status[2581] = `IFUPATH645.swl.thr1_state;
thread_status[2582] = `IFUPATH645.swl.thr2_state;
thread_status[2583] = `IFUPATH645.swl.thr3_state;
thread_status[2584] = `IFUPATH646.swl.thr0_state;
thread_status[2585] = `IFUPATH646.swl.thr1_state;
thread_status[2586] = `IFUPATH646.swl.thr2_state;
thread_status[2587] = `IFUPATH646.swl.thr3_state;
thread_status[2588] = `IFUPATH647.swl.thr0_state;
thread_status[2589] = `IFUPATH647.swl.thr1_state;
thread_status[2590] = `IFUPATH647.swl.thr2_state;
thread_status[2591] = `IFUPATH647.swl.thr3_state;
thread_status[2592] = `IFUPATH648.swl.thr0_state;
thread_status[2593] = `IFUPATH648.swl.thr1_state;
thread_status[2594] = `IFUPATH648.swl.thr2_state;
thread_status[2595] = `IFUPATH648.swl.thr3_state;
thread_status[2596] = `IFUPATH649.swl.thr0_state;
thread_status[2597] = `IFUPATH649.swl.thr1_state;
thread_status[2598] = `IFUPATH649.swl.thr2_state;
thread_status[2599] = `IFUPATH649.swl.thr3_state;
thread_status[2600] = `IFUPATH650.swl.thr0_state;
thread_status[2601] = `IFUPATH650.swl.thr1_state;
thread_status[2602] = `IFUPATH650.swl.thr2_state;
thread_status[2603] = `IFUPATH650.swl.thr3_state;
thread_status[2604] = `IFUPATH651.swl.thr0_state;
thread_status[2605] = `IFUPATH651.swl.thr1_state;
thread_status[2606] = `IFUPATH651.swl.thr2_state;
thread_status[2607] = `IFUPATH651.swl.thr3_state;
thread_status[2608] = `IFUPATH652.swl.thr0_state;
thread_status[2609] = `IFUPATH652.swl.thr1_state;
thread_status[2610] = `IFUPATH652.swl.thr2_state;
thread_status[2611] = `IFUPATH652.swl.thr3_state;
thread_status[2612] = `IFUPATH653.swl.thr0_state;
thread_status[2613] = `IFUPATH653.swl.thr1_state;
thread_status[2614] = `IFUPATH653.swl.thr2_state;
thread_status[2615] = `IFUPATH653.swl.thr3_state;
thread_status[2616] = `IFUPATH654.swl.thr0_state;
thread_status[2617] = `IFUPATH654.swl.thr1_state;
thread_status[2618] = `IFUPATH654.swl.thr2_state;
thread_status[2619] = `IFUPATH654.swl.thr3_state;
thread_status[2620] = `IFUPATH655.swl.thr0_state;
thread_status[2621] = `IFUPATH655.swl.thr1_state;
thread_status[2622] = `IFUPATH655.swl.thr2_state;
thread_status[2623] = `IFUPATH655.swl.thr3_state;
thread_status[2624] = `IFUPATH656.swl.thr0_state;
thread_status[2625] = `IFUPATH656.swl.thr1_state;
thread_status[2626] = `IFUPATH656.swl.thr2_state;
thread_status[2627] = `IFUPATH656.swl.thr3_state;
thread_status[2628] = `IFUPATH657.swl.thr0_state;
thread_status[2629] = `IFUPATH657.swl.thr1_state;
thread_status[2630] = `IFUPATH657.swl.thr2_state;
thread_status[2631] = `IFUPATH657.swl.thr3_state;
thread_status[2632] = `IFUPATH658.swl.thr0_state;
thread_status[2633] = `IFUPATH658.swl.thr1_state;
thread_status[2634] = `IFUPATH658.swl.thr2_state;
thread_status[2635] = `IFUPATH658.swl.thr3_state;
thread_status[2636] = `IFUPATH659.swl.thr0_state;
thread_status[2637] = `IFUPATH659.swl.thr1_state;
thread_status[2638] = `IFUPATH659.swl.thr2_state;
thread_status[2639] = `IFUPATH659.swl.thr3_state;
thread_status[2640] = `IFUPATH660.swl.thr0_state;
thread_status[2641] = `IFUPATH660.swl.thr1_state;
thread_status[2642] = `IFUPATH660.swl.thr2_state;
thread_status[2643] = `IFUPATH660.swl.thr3_state;
thread_status[2644] = `IFUPATH661.swl.thr0_state;
thread_status[2645] = `IFUPATH661.swl.thr1_state;
thread_status[2646] = `IFUPATH661.swl.thr2_state;
thread_status[2647] = `IFUPATH661.swl.thr3_state;
thread_status[2648] = `IFUPATH662.swl.thr0_state;
thread_status[2649] = `IFUPATH662.swl.thr1_state;
thread_status[2650] = `IFUPATH662.swl.thr2_state;
thread_status[2651] = `IFUPATH662.swl.thr3_state;
thread_status[2652] = `IFUPATH663.swl.thr0_state;
thread_status[2653] = `IFUPATH663.swl.thr1_state;
thread_status[2654] = `IFUPATH663.swl.thr2_state;
thread_status[2655] = `IFUPATH663.swl.thr3_state;
thread_status[2656] = `IFUPATH664.swl.thr0_state;
thread_status[2657] = `IFUPATH664.swl.thr1_state;
thread_status[2658] = `IFUPATH664.swl.thr2_state;
thread_status[2659] = `IFUPATH664.swl.thr3_state;
thread_status[2660] = `IFUPATH665.swl.thr0_state;
thread_status[2661] = `IFUPATH665.swl.thr1_state;
thread_status[2662] = `IFUPATH665.swl.thr2_state;
thread_status[2663] = `IFUPATH665.swl.thr3_state;
thread_status[2664] = `IFUPATH666.swl.thr0_state;
thread_status[2665] = `IFUPATH666.swl.thr1_state;
thread_status[2666] = `IFUPATH666.swl.thr2_state;
thread_status[2667] = `IFUPATH666.swl.thr3_state;
thread_status[2668] = `IFUPATH667.swl.thr0_state;
thread_status[2669] = `IFUPATH667.swl.thr1_state;
thread_status[2670] = `IFUPATH667.swl.thr2_state;
thread_status[2671] = `IFUPATH667.swl.thr3_state;
thread_status[2672] = `IFUPATH668.swl.thr0_state;
thread_status[2673] = `IFUPATH668.swl.thr1_state;
thread_status[2674] = `IFUPATH668.swl.thr2_state;
thread_status[2675] = `IFUPATH668.swl.thr3_state;
thread_status[2676] = `IFUPATH669.swl.thr0_state;
thread_status[2677] = `IFUPATH669.swl.thr1_state;
thread_status[2678] = `IFUPATH669.swl.thr2_state;
thread_status[2679] = `IFUPATH669.swl.thr3_state;
thread_status[2680] = `IFUPATH670.swl.thr0_state;
thread_status[2681] = `IFUPATH670.swl.thr1_state;
thread_status[2682] = `IFUPATH670.swl.thr2_state;
thread_status[2683] = `IFUPATH670.swl.thr3_state;
thread_status[2684] = `IFUPATH671.swl.thr0_state;
thread_status[2685] = `IFUPATH671.swl.thr1_state;
thread_status[2686] = `IFUPATH671.swl.thr2_state;
thread_status[2687] = `IFUPATH671.swl.thr3_state;
thread_status[2688] = `IFUPATH672.swl.thr0_state;
thread_status[2689] = `IFUPATH672.swl.thr1_state;
thread_status[2690] = `IFUPATH672.swl.thr2_state;
thread_status[2691] = `IFUPATH672.swl.thr3_state;
thread_status[2692] = `IFUPATH673.swl.thr0_state;
thread_status[2693] = `IFUPATH673.swl.thr1_state;
thread_status[2694] = `IFUPATH673.swl.thr2_state;
thread_status[2695] = `IFUPATH673.swl.thr3_state;
thread_status[2696] = `IFUPATH674.swl.thr0_state;
thread_status[2697] = `IFUPATH674.swl.thr1_state;
thread_status[2698] = `IFUPATH674.swl.thr2_state;
thread_status[2699] = `IFUPATH674.swl.thr3_state;
thread_status[2700] = `IFUPATH675.swl.thr0_state;
thread_status[2701] = `IFUPATH675.swl.thr1_state;
thread_status[2702] = `IFUPATH675.swl.thr2_state;
thread_status[2703] = `IFUPATH675.swl.thr3_state;
thread_status[2704] = `IFUPATH676.swl.thr0_state;
thread_status[2705] = `IFUPATH676.swl.thr1_state;
thread_status[2706] = `IFUPATH676.swl.thr2_state;
thread_status[2707] = `IFUPATH676.swl.thr3_state;
thread_status[2708] = `IFUPATH677.swl.thr0_state;
thread_status[2709] = `IFUPATH677.swl.thr1_state;
thread_status[2710] = `IFUPATH677.swl.thr2_state;
thread_status[2711] = `IFUPATH677.swl.thr3_state;
thread_status[2712] = `IFUPATH678.swl.thr0_state;
thread_status[2713] = `IFUPATH678.swl.thr1_state;
thread_status[2714] = `IFUPATH678.swl.thr2_state;
thread_status[2715] = `IFUPATH678.swl.thr3_state;
thread_status[2716] = `IFUPATH679.swl.thr0_state;
thread_status[2717] = `IFUPATH679.swl.thr1_state;
thread_status[2718] = `IFUPATH679.swl.thr2_state;
thread_status[2719] = `IFUPATH679.swl.thr3_state;
thread_status[2720] = `IFUPATH680.swl.thr0_state;
thread_status[2721] = `IFUPATH680.swl.thr1_state;
thread_status[2722] = `IFUPATH680.swl.thr2_state;
thread_status[2723] = `IFUPATH680.swl.thr3_state;
thread_status[2724] = `IFUPATH681.swl.thr0_state;
thread_status[2725] = `IFUPATH681.swl.thr1_state;
thread_status[2726] = `IFUPATH681.swl.thr2_state;
thread_status[2727] = `IFUPATH681.swl.thr3_state;
thread_status[2728] = `IFUPATH682.swl.thr0_state;
thread_status[2729] = `IFUPATH682.swl.thr1_state;
thread_status[2730] = `IFUPATH682.swl.thr2_state;
thread_status[2731] = `IFUPATH682.swl.thr3_state;
thread_status[2732] = `IFUPATH683.swl.thr0_state;
thread_status[2733] = `IFUPATH683.swl.thr1_state;
thread_status[2734] = `IFUPATH683.swl.thr2_state;
thread_status[2735] = `IFUPATH683.swl.thr3_state;
thread_status[2736] = `IFUPATH684.swl.thr0_state;
thread_status[2737] = `IFUPATH684.swl.thr1_state;
thread_status[2738] = `IFUPATH684.swl.thr2_state;
thread_status[2739] = `IFUPATH684.swl.thr3_state;
thread_status[2740] = `IFUPATH685.swl.thr0_state;
thread_status[2741] = `IFUPATH685.swl.thr1_state;
thread_status[2742] = `IFUPATH685.swl.thr2_state;
thread_status[2743] = `IFUPATH685.swl.thr3_state;
thread_status[2744] = `IFUPATH686.swl.thr0_state;
thread_status[2745] = `IFUPATH686.swl.thr1_state;
thread_status[2746] = `IFUPATH686.swl.thr2_state;
thread_status[2747] = `IFUPATH686.swl.thr3_state;
thread_status[2748] = `IFUPATH687.swl.thr0_state;
thread_status[2749] = `IFUPATH687.swl.thr1_state;
thread_status[2750] = `IFUPATH687.swl.thr2_state;
thread_status[2751] = `IFUPATH687.swl.thr3_state;
thread_status[2752] = `IFUPATH688.swl.thr0_state;
thread_status[2753] = `IFUPATH688.swl.thr1_state;
thread_status[2754] = `IFUPATH688.swl.thr2_state;
thread_status[2755] = `IFUPATH688.swl.thr3_state;
thread_status[2756] = `IFUPATH689.swl.thr0_state;
thread_status[2757] = `IFUPATH689.swl.thr1_state;
thread_status[2758] = `IFUPATH689.swl.thr2_state;
thread_status[2759] = `IFUPATH689.swl.thr3_state;
thread_status[2760] = `IFUPATH690.swl.thr0_state;
thread_status[2761] = `IFUPATH690.swl.thr1_state;
thread_status[2762] = `IFUPATH690.swl.thr2_state;
thread_status[2763] = `IFUPATH690.swl.thr3_state;
thread_status[2764] = `IFUPATH691.swl.thr0_state;
thread_status[2765] = `IFUPATH691.swl.thr1_state;
thread_status[2766] = `IFUPATH691.swl.thr2_state;
thread_status[2767] = `IFUPATH691.swl.thr3_state;
thread_status[2768] = `IFUPATH692.swl.thr0_state;
thread_status[2769] = `IFUPATH692.swl.thr1_state;
thread_status[2770] = `IFUPATH692.swl.thr2_state;
thread_status[2771] = `IFUPATH692.swl.thr3_state;
thread_status[2772] = `IFUPATH693.swl.thr0_state;
thread_status[2773] = `IFUPATH693.swl.thr1_state;
thread_status[2774] = `IFUPATH693.swl.thr2_state;
thread_status[2775] = `IFUPATH693.swl.thr3_state;
thread_status[2776] = `IFUPATH694.swl.thr0_state;
thread_status[2777] = `IFUPATH694.swl.thr1_state;
thread_status[2778] = `IFUPATH694.swl.thr2_state;
thread_status[2779] = `IFUPATH694.swl.thr3_state;
thread_status[2780] = `IFUPATH695.swl.thr0_state;
thread_status[2781] = `IFUPATH695.swl.thr1_state;
thread_status[2782] = `IFUPATH695.swl.thr2_state;
thread_status[2783] = `IFUPATH695.swl.thr3_state;
thread_status[2784] = `IFUPATH696.swl.thr0_state;
thread_status[2785] = `IFUPATH696.swl.thr1_state;
thread_status[2786] = `IFUPATH696.swl.thr2_state;
thread_status[2787] = `IFUPATH696.swl.thr3_state;
thread_status[2788] = `IFUPATH697.swl.thr0_state;
thread_status[2789] = `IFUPATH697.swl.thr1_state;
thread_status[2790] = `IFUPATH697.swl.thr2_state;
thread_status[2791] = `IFUPATH697.swl.thr3_state;
thread_status[2792] = `IFUPATH698.swl.thr0_state;
thread_status[2793] = `IFUPATH698.swl.thr1_state;
thread_status[2794] = `IFUPATH698.swl.thr2_state;
thread_status[2795] = `IFUPATH698.swl.thr3_state;
thread_status[2796] = `IFUPATH699.swl.thr0_state;
thread_status[2797] = `IFUPATH699.swl.thr1_state;
thread_status[2798] = `IFUPATH699.swl.thr2_state;
thread_status[2799] = `IFUPATH699.swl.thr3_state;
thread_status[2800] = `IFUPATH700.swl.thr0_state;
thread_status[2801] = `IFUPATH700.swl.thr1_state;
thread_status[2802] = `IFUPATH700.swl.thr2_state;
thread_status[2803] = `IFUPATH700.swl.thr3_state;
thread_status[2804] = `IFUPATH701.swl.thr0_state;
thread_status[2805] = `IFUPATH701.swl.thr1_state;
thread_status[2806] = `IFUPATH701.swl.thr2_state;
thread_status[2807] = `IFUPATH701.swl.thr3_state;
thread_status[2808] = `IFUPATH702.swl.thr0_state;
thread_status[2809] = `IFUPATH702.swl.thr1_state;
thread_status[2810] = `IFUPATH702.swl.thr2_state;
thread_status[2811] = `IFUPATH702.swl.thr3_state;
thread_status[2812] = `IFUPATH703.swl.thr0_state;
thread_status[2813] = `IFUPATH703.swl.thr1_state;
thread_status[2814] = `IFUPATH703.swl.thr2_state;
thread_status[2815] = `IFUPATH703.swl.thr3_state;
thread_status[2816] = `IFUPATH704.swl.thr0_state;
thread_status[2817] = `IFUPATH704.swl.thr1_state;
thread_status[2818] = `IFUPATH704.swl.thr2_state;
thread_status[2819] = `IFUPATH704.swl.thr3_state;
thread_status[2820] = `IFUPATH705.swl.thr0_state;
thread_status[2821] = `IFUPATH705.swl.thr1_state;
thread_status[2822] = `IFUPATH705.swl.thr2_state;
thread_status[2823] = `IFUPATH705.swl.thr3_state;
thread_status[2824] = `IFUPATH706.swl.thr0_state;
thread_status[2825] = `IFUPATH706.swl.thr1_state;
thread_status[2826] = `IFUPATH706.swl.thr2_state;
thread_status[2827] = `IFUPATH706.swl.thr3_state;
thread_status[2828] = `IFUPATH707.swl.thr0_state;
thread_status[2829] = `IFUPATH707.swl.thr1_state;
thread_status[2830] = `IFUPATH707.swl.thr2_state;
thread_status[2831] = `IFUPATH707.swl.thr3_state;
thread_status[2832] = `IFUPATH708.swl.thr0_state;
thread_status[2833] = `IFUPATH708.swl.thr1_state;
thread_status[2834] = `IFUPATH708.swl.thr2_state;
thread_status[2835] = `IFUPATH708.swl.thr3_state;
thread_status[2836] = `IFUPATH709.swl.thr0_state;
thread_status[2837] = `IFUPATH709.swl.thr1_state;
thread_status[2838] = `IFUPATH709.swl.thr2_state;
thread_status[2839] = `IFUPATH709.swl.thr3_state;
thread_status[2840] = `IFUPATH710.swl.thr0_state;
thread_status[2841] = `IFUPATH710.swl.thr1_state;
thread_status[2842] = `IFUPATH710.swl.thr2_state;
thread_status[2843] = `IFUPATH710.swl.thr3_state;
thread_status[2844] = `IFUPATH711.swl.thr0_state;
thread_status[2845] = `IFUPATH711.swl.thr1_state;
thread_status[2846] = `IFUPATH711.swl.thr2_state;
thread_status[2847] = `IFUPATH711.swl.thr3_state;
thread_status[2848] = `IFUPATH712.swl.thr0_state;
thread_status[2849] = `IFUPATH712.swl.thr1_state;
thread_status[2850] = `IFUPATH712.swl.thr2_state;
thread_status[2851] = `IFUPATH712.swl.thr3_state;
thread_status[2852] = `IFUPATH713.swl.thr0_state;
thread_status[2853] = `IFUPATH713.swl.thr1_state;
thread_status[2854] = `IFUPATH713.swl.thr2_state;
thread_status[2855] = `IFUPATH713.swl.thr3_state;
thread_status[2856] = `IFUPATH714.swl.thr0_state;
thread_status[2857] = `IFUPATH714.swl.thr1_state;
thread_status[2858] = `IFUPATH714.swl.thr2_state;
thread_status[2859] = `IFUPATH714.swl.thr3_state;
thread_status[2860] = `IFUPATH715.swl.thr0_state;
thread_status[2861] = `IFUPATH715.swl.thr1_state;
thread_status[2862] = `IFUPATH715.swl.thr2_state;
thread_status[2863] = `IFUPATH715.swl.thr3_state;
thread_status[2864] = `IFUPATH716.swl.thr0_state;
thread_status[2865] = `IFUPATH716.swl.thr1_state;
thread_status[2866] = `IFUPATH716.swl.thr2_state;
thread_status[2867] = `IFUPATH716.swl.thr3_state;
thread_status[2868] = `IFUPATH717.swl.thr0_state;
thread_status[2869] = `IFUPATH717.swl.thr1_state;
thread_status[2870] = `IFUPATH717.swl.thr2_state;
thread_status[2871] = `IFUPATH717.swl.thr3_state;
thread_status[2872] = `IFUPATH718.swl.thr0_state;
thread_status[2873] = `IFUPATH718.swl.thr1_state;
thread_status[2874] = `IFUPATH718.swl.thr2_state;
thread_status[2875] = `IFUPATH718.swl.thr3_state;
thread_status[2876] = `IFUPATH719.swl.thr0_state;
thread_status[2877] = `IFUPATH719.swl.thr1_state;
thread_status[2878] = `IFUPATH719.swl.thr2_state;
thread_status[2879] = `IFUPATH719.swl.thr3_state;
thread_status[2880] = `IFUPATH720.swl.thr0_state;
thread_status[2881] = `IFUPATH720.swl.thr1_state;
thread_status[2882] = `IFUPATH720.swl.thr2_state;
thread_status[2883] = `IFUPATH720.swl.thr3_state;
thread_status[2884] = `IFUPATH721.swl.thr0_state;
thread_status[2885] = `IFUPATH721.swl.thr1_state;
thread_status[2886] = `IFUPATH721.swl.thr2_state;
thread_status[2887] = `IFUPATH721.swl.thr3_state;
thread_status[2888] = `IFUPATH722.swl.thr0_state;
thread_status[2889] = `IFUPATH722.swl.thr1_state;
thread_status[2890] = `IFUPATH722.swl.thr2_state;
thread_status[2891] = `IFUPATH722.swl.thr3_state;
thread_status[2892] = `IFUPATH723.swl.thr0_state;
thread_status[2893] = `IFUPATH723.swl.thr1_state;
thread_status[2894] = `IFUPATH723.swl.thr2_state;
thread_status[2895] = `IFUPATH723.swl.thr3_state;
thread_status[2896] = `IFUPATH724.swl.thr0_state;
thread_status[2897] = `IFUPATH724.swl.thr1_state;
thread_status[2898] = `IFUPATH724.swl.thr2_state;
thread_status[2899] = `IFUPATH724.swl.thr3_state;
thread_status[2900] = `IFUPATH725.swl.thr0_state;
thread_status[2901] = `IFUPATH725.swl.thr1_state;
thread_status[2902] = `IFUPATH725.swl.thr2_state;
thread_status[2903] = `IFUPATH725.swl.thr3_state;
thread_status[2904] = `IFUPATH726.swl.thr0_state;
thread_status[2905] = `IFUPATH726.swl.thr1_state;
thread_status[2906] = `IFUPATH726.swl.thr2_state;
thread_status[2907] = `IFUPATH726.swl.thr3_state;
thread_status[2908] = `IFUPATH727.swl.thr0_state;
thread_status[2909] = `IFUPATH727.swl.thr1_state;
thread_status[2910] = `IFUPATH727.swl.thr2_state;
thread_status[2911] = `IFUPATH727.swl.thr3_state;
thread_status[2912] = `IFUPATH728.swl.thr0_state;
thread_status[2913] = `IFUPATH728.swl.thr1_state;
thread_status[2914] = `IFUPATH728.swl.thr2_state;
thread_status[2915] = `IFUPATH728.swl.thr3_state;
thread_status[2916] = `IFUPATH729.swl.thr0_state;
thread_status[2917] = `IFUPATH729.swl.thr1_state;
thread_status[2918] = `IFUPATH729.swl.thr2_state;
thread_status[2919] = `IFUPATH729.swl.thr3_state;
thread_status[2920] = `IFUPATH730.swl.thr0_state;
thread_status[2921] = `IFUPATH730.swl.thr1_state;
thread_status[2922] = `IFUPATH730.swl.thr2_state;
thread_status[2923] = `IFUPATH730.swl.thr3_state;
thread_status[2924] = `IFUPATH731.swl.thr0_state;
thread_status[2925] = `IFUPATH731.swl.thr1_state;
thread_status[2926] = `IFUPATH731.swl.thr2_state;
thread_status[2927] = `IFUPATH731.swl.thr3_state;
thread_status[2928] = `IFUPATH732.swl.thr0_state;
thread_status[2929] = `IFUPATH732.swl.thr1_state;
thread_status[2930] = `IFUPATH732.swl.thr2_state;
thread_status[2931] = `IFUPATH732.swl.thr3_state;
thread_status[2932] = `IFUPATH733.swl.thr0_state;
thread_status[2933] = `IFUPATH733.swl.thr1_state;
thread_status[2934] = `IFUPATH733.swl.thr2_state;
thread_status[2935] = `IFUPATH733.swl.thr3_state;
thread_status[2936] = `IFUPATH734.swl.thr0_state;
thread_status[2937] = `IFUPATH734.swl.thr1_state;
thread_status[2938] = `IFUPATH734.swl.thr2_state;
thread_status[2939] = `IFUPATH734.swl.thr3_state;
thread_status[2940] = `IFUPATH735.swl.thr0_state;
thread_status[2941] = `IFUPATH735.swl.thr1_state;
thread_status[2942] = `IFUPATH735.swl.thr2_state;
thread_status[2943] = `IFUPATH735.swl.thr3_state;
thread_status[2944] = `IFUPATH736.swl.thr0_state;
thread_status[2945] = `IFUPATH736.swl.thr1_state;
thread_status[2946] = `IFUPATH736.swl.thr2_state;
thread_status[2947] = `IFUPATH736.swl.thr3_state;
thread_status[2948] = `IFUPATH737.swl.thr0_state;
thread_status[2949] = `IFUPATH737.swl.thr1_state;
thread_status[2950] = `IFUPATH737.swl.thr2_state;
thread_status[2951] = `IFUPATH737.swl.thr3_state;
thread_status[2952] = `IFUPATH738.swl.thr0_state;
thread_status[2953] = `IFUPATH738.swl.thr1_state;
thread_status[2954] = `IFUPATH738.swl.thr2_state;
thread_status[2955] = `IFUPATH738.swl.thr3_state;
thread_status[2956] = `IFUPATH739.swl.thr0_state;
thread_status[2957] = `IFUPATH739.swl.thr1_state;
thread_status[2958] = `IFUPATH739.swl.thr2_state;
thread_status[2959] = `IFUPATH739.swl.thr3_state;
thread_status[2960] = `IFUPATH740.swl.thr0_state;
thread_status[2961] = `IFUPATH740.swl.thr1_state;
thread_status[2962] = `IFUPATH740.swl.thr2_state;
thread_status[2963] = `IFUPATH740.swl.thr3_state;
thread_status[2964] = `IFUPATH741.swl.thr0_state;
thread_status[2965] = `IFUPATH741.swl.thr1_state;
thread_status[2966] = `IFUPATH741.swl.thr2_state;
thread_status[2967] = `IFUPATH741.swl.thr3_state;
thread_status[2968] = `IFUPATH742.swl.thr0_state;
thread_status[2969] = `IFUPATH742.swl.thr1_state;
thread_status[2970] = `IFUPATH742.swl.thr2_state;
thread_status[2971] = `IFUPATH742.swl.thr3_state;
thread_status[2972] = `IFUPATH743.swl.thr0_state;
thread_status[2973] = `IFUPATH743.swl.thr1_state;
thread_status[2974] = `IFUPATH743.swl.thr2_state;
thread_status[2975] = `IFUPATH743.swl.thr3_state;
thread_status[2976] = `IFUPATH744.swl.thr0_state;
thread_status[2977] = `IFUPATH744.swl.thr1_state;
thread_status[2978] = `IFUPATH744.swl.thr2_state;
thread_status[2979] = `IFUPATH744.swl.thr3_state;
thread_status[2980] = `IFUPATH745.swl.thr0_state;
thread_status[2981] = `IFUPATH745.swl.thr1_state;
thread_status[2982] = `IFUPATH745.swl.thr2_state;
thread_status[2983] = `IFUPATH745.swl.thr3_state;
thread_status[2984] = `IFUPATH746.swl.thr0_state;
thread_status[2985] = `IFUPATH746.swl.thr1_state;
thread_status[2986] = `IFUPATH746.swl.thr2_state;
thread_status[2987] = `IFUPATH746.swl.thr3_state;
thread_status[2988] = `IFUPATH747.swl.thr0_state;
thread_status[2989] = `IFUPATH747.swl.thr1_state;
thread_status[2990] = `IFUPATH747.swl.thr2_state;
thread_status[2991] = `IFUPATH747.swl.thr3_state;
thread_status[2992] = `IFUPATH748.swl.thr0_state;
thread_status[2993] = `IFUPATH748.swl.thr1_state;
thread_status[2994] = `IFUPATH748.swl.thr2_state;
thread_status[2995] = `IFUPATH748.swl.thr3_state;
thread_status[2996] = `IFUPATH749.swl.thr0_state;
thread_status[2997] = `IFUPATH749.swl.thr1_state;
thread_status[2998] = `IFUPATH749.swl.thr2_state;
thread_status[2999] = `IFUPATH749.swl.thr3_state;
thread_status[3000] = `IFUPATH750.swl.thr0_state;
thread_status[3001] = `IFUPATH750.swl.thr1_state;
thread_status[3002] = `IFUPATH750.swl.thr2_state;
thread_status[3003] = `IFUPATH750.swl.thr3_state;
thread_status[3004] = `IFUPATH751.swl.thr0_state;
thread_status[3005] = `IFUPATH751.swl.thr1_state;
thread_status[3006] = `IFUPATH751.swl.thr2_state;
thread_status[3007] = `IFUPATH751.swl.thr3_state;
thread_status[3008] = `IFUPATH752.swl.thr0_state;
thread_status[3009] = `IFUPATH752.swl.thr1_state;
thread_status[3010] = `IFUPATH752.swl.thr2_state;
thread_status[3011] = `IFUPATH752.swl.thr3_state;
thread_status[3012] = `IFUPATH753.swl.thr0_state;
thread_status[3013] = `IFUPATH753.swl.thr1_state;
thread_status[3014] = `IFUPATH753.swl.thr2_state;
thread_status[3015] = `IFUPATH753.swl.thr3_state;
thread_status[3016] = `IFUPATH754.swl.thr0_state;
thread_status[3017] = `IFUPATH754.swl.thr1_state;
thread_status[3018] = `IFUPATH754.swl.thr2_state;
thread_status[3019] = `IFUPATH754.swl.thr3_state;
thread_status[3020] = `IFUPATH755.swl.thr0_state;
thread_status[3021] = `IFUPATH755.swl.thr1_state;
thread_status[3022] = `IFUPATH755.swl.thr2_state;
thread_status[3023] = `IFUPATH755.swl.thr3_state;
thread_status[3024] = `IFUPATH756.swl.thr0_state;
thread_status[3025] = `IFUPATH756.swl.thr1_state;
thread_status[3026] = `IFUPATH756.swl.thr2_state;
thread_status[3027] = `IFUPATH756.swl.thr3_state;
thread_status[3028] = `IFUPATH757.swl.thr0_state;
thread_status[3029] = `IFUPATH757.swl.thr1_state;
thread_status[3030] = `IFUPATH757.swl.thr2_state;
thread_status[3031] = `IFUPATH757.swl.thr3_state;
thread_status[3032] = `IFUPATH758.swl.thr0_state;
thread_status[3033] = `IFUPATH758.swl.thr1_state;
thread_status[3034] = `IFUPATH758.swl.thr2_state;
thread_status[3035] = `IFUPATH758.swl.thr3_state;
thread_status[3036] = `IFUPATH759.swl.thr0_state;
thread_status[3037] = `IFUPATH759.swl.thr1_state;
thread_status[3038] = `IFUPATH759.swl.thr2_state;
thread_status[3039] = `IFUPATH759.swl.thr3_state;
thread_status[3040] = `IFUPATH760.swl.thr0_state;
thread_status[3041] = `IFUPATH760.swl.thr1_state;
thread_status[3042] = `IFUPATH760.swl.thr2_state;
thread_status[3043] = `IFUPATH760.swl.thr3_state;
thread_status[3044] = `IFUPATH761.swl.thr0_state;
thread_status[3045] = `IFUPATH761.swl.thr1_state;
thread_status[3046] = `IFUPATH761.swl.thr2_state;
thread_status[3047] = `IFUPATH761.swl.thr3_state;
thread_status[3048] = `IFUPATH762.swl.thr0_state;
thread_status[3049] = `IFUPATH762.swl.thr1_state;
thread_status[3050] = `IFUPATH762.swl.thr2_state;
thread_status[3051] = `IFUPATH762.swl.thr3_state;
thread_status[3052] = `IFUPATH763.swl.thr0_state;
thread_status[3053] = `IFUPATH763.swl.thr1_state;
thread_status[3054] = `IFUPATH763.swl.thr2_state;
thread_status[3055] = `IFUPATH763.swl.thr3_state;
thread_status[3056] = `IFUPATH764.swl.thr0_state;
thread_status[3057] = `IFUPATH764.swl.thr1_state;
thread_status[3058] = `IFUPATH764.swl.thr2_state;
thread_status[3059] = `IFUPATH764.swl.thr3_state;
thread_status[3060] = `IFUPATH765.swl.thr0_state;
thread_status[3061] = `IFUPATH765.swl.thr1_state;
thread_status[3062] = `IFUPATH765.swl.thr2_state;
thread_status[3063] = `IFUPATH765.swl.thr3_state;
thread_status[3064] = `IFUPATH766.swl.thr0_state;
thread_status[3065] = `IFUPATH766.swl.thr1_state;
thread_status[3066] = `IFUPATH766.swl.thr2_state;
thread_status[3067] = `IFUPATH766.swl.thr3_state;
thread_status[3068] = `IFUPATH767.swl.thr0_state;
thread_status[3069] = `IFUPATH767.swl.thr1_state;
thread_status[3070] = `IFUPATH767.swl.thr2_state;
thread_status[3071] = `IFUPATH767.swl.thr3_state;
thread_status[3072] = `IFUPATH768.swl.thr0_state;
thread_status[3073] = `IFUPATH768.swl.thr1_state;
thread_status[3074] = `IFUPATH768.swl.thr2_state;
thread_status[3075] = `IFUPATH768.swl.thr3_state;
thread_status[3076] = `IFUPATH769.swl.thr0_state;
thread_status[3077] = `IFUPATH769.swl.thr1_state;
thread_status[3078] = `IFUPATH769.swl.thr2_state;
thread_status[3079] = `IFUPATH769.swl.thr3_state;
thread_status[3080] = `IFUPATH770.swl.thr0_state;
thread_status[3081] = `IFUPATH770.swl.thr1_state;
thread_status[3082] = `IFUPATH770.swl.thr2_state;
thread_status[3083] = `IFUPATH770.swl.thr3_state;
thread_status[3084] = `IFUPATH771.swl.thr0_state;
thread_status[3085] = `IFUPATH771.swl.thr1_state;
thread_status[3086] = `IFUPATH771.swl.thr2_state;
thread_status[3087] = `IFUPATH771.swl.thr3_state;
thread_status[3088] = `IFUPATH772.swl.thr0_state;
thread_status[3089] = `IFUPATH772.swl.thr1_state;
thread_status[3090] = `IFUPATH772.swl.thr2_state;
thread_status[3091] = `IFUPATH772.swl.thr3_state;
thread_status[3092] = `IFUPATH773.swl.thr0_state;
thread_status[3093] = `IFUPATH773.swl.thr1_state;
thread_status[3094] = `IFUPATH773.swl.thr2_state;
thread_status[3095] = `IFUPATH773.swl.thr3_state;
thread_status[3096] = `IFUPATH774.swl.thr0_state;
thread_status[3097] = `IFUPATH774.swl.thr1_state;
thread_status[3098] = `IFUPATH774.swl.thr2_state;
thread_status[3099] = `IFUPATH774.swl.thr3_state;
thread_status[3100] = `IFUPATH775.swl.thr0_state;
thread_status[3101] = `IFUPATH775.swl.thr1_state;
thread_status[3102] = `IFUPATH775.swl.thr2_state;
thread_status[3103] = `IFUPATH775.swl.thr3_state;
thread_status[3104] = `IFUPATH776.swl.thr0_state;
thread_status[3105] = `IFUPATH776.swl.thr1_state;
thread_status[3106] = `IFUPATH776.swl.thr2_state;
thread_status[3107] = `IFUPATH776.swl.thr3_state;
thread_status[3108] = `IFUPATH777.swl.thr0_state;
thread_status[3109] = `IFUPATH777.swl.thr1_state;
thread_status[3110] = `IFUPATH777.swl.thr2_state;
thread_status[3111] = `IFUPATH777.swl.thr3_state;
thread_status[3112] = `IFUPATH778.swl.thr0_state;
thread_status[3113] = `IFUPATH778.swl.thr1_state;
thread_status[3114] = `IFUPATH778.swl.thr2_state;
thread_status[3115] = `IFUPATH778.swl.thr3_state;
thread_status[3116] = `IFUPATH779.swl.thr0_state;
thread_status[3117] = `IFUPATH779.swl.thr1_state;
thread_status[3118] = `IFUPATH779.swl.thr2_state;
thread_status[3119] = `IFUPATH779.swl.thr3_state;
thread_status[3120] = `IFUPATH780.swl.thr0_state;
thread_status[3121] = `IFUPATH780.swl.thr1_state;
thread_status[3122] = `IFUPATH780.swl.thr2_state;
thread_status[3123] = `IFUPATH780.swl.thr3_state;
thread_status[3124] = `IFUPATH781.swl.thr0_state;
thread_status[3125] = `IFUPATH781.swl.thr1_state;
thread_status[3126] = `IFUPATH781.swl.thr2_state;
thread_status[3127] = `IFUPATH781.swl.thr3_state;
thread_status[3128] = `IFUPATH782.swl.thr0_state;
thread_status[3129] = `IFUPATH782.swl.thr1_state;
thread_status[3130] = `IFUPATH782.swl.thr2_state;
thread_status[3131] = `IFUPATH782.swl.thr3_state;
thread_status[3132] = `IFUPATH783.swl.thr0_state;
thread_status[3133] = `IFUPATH783.swl.thr1_state;
thread_status[3134] = `IFUPATH783.swl.thr2_state;
thread_status[3135] = `IFUPATH783.swl.thr3_state;
thread_status[3136] = `IFUPATH784.swl.thr0_state;
thread_status[3137] = `IFUPATH784.swl.thr1_state;
thread_status[3138] = `IFUPATH784.swl.thr2_state;
thread_status[3139] = `IFUPATH784.swl.thr3_state;
thread_status[3140] = `IFUPATH785.swl.thr0_state;
thread_status[3141] = `IFUPATH785.swl.thr1_state;
thread_status[3142] = `IFUPATH785.swl.thr2_state;
thread_status[3143] = `IFUPATH785.swl.thr3_state;
thread_status[3144] = `IFUPATH786.swl.thr0_state;
thread_status[3145] = `IFUPATH786.swl.thr1_state;
thread_status[3146] = `IFUPATH786.swl.thr2_state;
thread_status[3147] = `IFUPATH786.swl.thr3_state;
thread_status[3148] = `IFUPATH787.swl.thr0_state;
thread_status[3149] = `IFUPATH787.swl.thr1_state;
thread_status[3150] = `IFUPATH787.swl.thr2_state;
thread_status[3151] = `IFUPATH787.swl.thr3_state;
thread_status[3152] = `IFUPATH788.swl.thr0_state;
thread_status[3153] = `IFUPATH788.swl.thr1_state;
thread_status[3154] = `IFUPATH788.swl.thr2_state;
thread_status[3155] = `IFUPATH788.swl.thr3_state;
thread_status[3156] = `IFUPATH789.swl.thr0_state;
thread_status[3157] = `IFUPATH789.swl.thr1_state;
thread_status[3158] = `IFUPATH789.swl.thr2_state;
thread_status[3159] = `IFUPATH789.swl.thr3_state;
thread_status[3160] = `IFUPATH790.swl.thr0_state;
thread_status[3161] = `IFUPATH790.swl.thr1_state;
thread_status[3162] = `IFUPATH790.swl.thr2_state;
thread_status[3163] = `IFUPATH790.swl.thr3_state;
thread_status[3164] = `IFUPATH791.swl.thr0_state;
thread_status[3165] = `IFUPATH791.swl.thr1_state;
thread_status[3166] = `IFUPATH791.swl.thr2_state;
thread_status[3167] = `IFUPATH791.swl.thr3_state;
thread_status[3168] = `IFUPATH792.swl.thr0_state;
thread_status[3169] = `IFUPATH792.swl.thr1_state;
thread_status[3170] = `IFUPATH792.swl.thr2_state;
thread_status[3171] = `IFUPATH792.swl.thr3_state;
thread_status[3172] = `IFUPATH793.swl.thr0_state;
thread_status[3173] = `IFUPATH793.swl.thr1_state;
thread_status[3174] = `IFUPATH793.swl.thr2_state;
thread_status[3175] = `IFUPATH793.swl.thr3_state;
thread_status[3176] = `IFUPATH794.swl.thr0_state;
thread_status[3177] = `IFUPATH794.swl.thr1_state;
thread_status[3178] = `IFUPATH794.swl.thr2_state;
thread_status[3179] = `IFUPATH794.swl.thr3_state;
thread_status[3180] = `IFUPATH795.swl.thr0_state;
thread_status[3181] = `IFUPATH795.swl.thr1_state;
thread_status[3182] = `IFUPATH795.swl.thr2_state;
thread_status[3183] = `IFUPATH795.swl.thr3_state;
thread_status[3184] = `IFUPATH796.swl.thr0_state;
thread_status[3185] = `IFUPATH796.swl.thr1_state;
thread_status[3186] = `IFUPATH796.swl.thr2_state;
thread_status[3187] = `IFUPATH796.swl.thr3_state;
thread_status[3188] = `IFUPATH797.swl.thr0_state;
thread_status[3189] = `IFUPATH797.swl.thr1_state;
thread_status[3190] = `IFUPATH797.swl.thr2_state;
thread_status[3191] = `IFUPATH797.swl.thr3_state;
thread_status[3192] = `IFUPATH798.swl.thr0_state;
thread_status[3193] = `IFUPATH798.swl.thr1_state;
thread_status[3194] = `IFUPATH798.swl.thr2_state;
thread_status[3195] = `IFUPATH798.swl.thr3_state;
thread_status[3196] = `IFUPATH799.swl.thr0_state;
thread_status[3197] = `IFUPATH799.swl.thr1_state;
thread_status[3198] = `IFUPATH799.swl.thr2_state;
thread_status[3199] = `IFUPATH799.swl.thr3_state;
thread_status[3200] = `IFUPATH800.swl.thr0_state;
thread_status[3201] = `IFUPATH800.swl.thr1_state;
thread_status[3202] = `IFUPATH800.swl.thr2_state;
thread_status[3203] = `IFUPATH800.swl.thr3_state;
thread_status[3204] = `IFUPATH801.swl.thr0_state;
thread_status[3205] = `IFUPATH801.swl.thr1_state;
thread_status[3206] = `IFUPATH801.swl.thr2_state;
thread_status[3207] = `IFUPATH801.swl.thr3_state;
thread_status[3208] = `IFUPATH802.swl.thr0_state;
thread_status[3209] = `IFUPATH802.swl.thr1_state;
thread_status[3210] = `IFUPATH802.swl.thr2_state;
thread_status[3211] = `IFUPATH802.swl.thr3_state;
thread_status[3212] = `IFUPATH803.swl.thr0_state;
thread_status[3213] = `IFUPATH803.swl.thr1_state;
thread_status[3214] = `IFUPATH803.swl.thr2_state;
thread_status[3215] = `IFUPATH803.swl.thr3_state;
thread_status[3216] = `IFUPATH804.swl.thr0_state;
thread_status[3217] = `IFUPATH804.swl.thr1_state;
thread_status[3218] = `IFUPATH804.swl.thr2_state;
thread_status[3219] = `IFUPATH804.swl.thr3_state;
thread_status[3220] = `IFUPATH805.swl.thr0_state;
thread_status[3221] = `IFUPATH805.swl.thr1_state;
thread_status[3222] = `IFUPATH805.swl.thr2_state;
thread_status[3223] = `IFUPATH805.swl.thr3_state;
thread_status[3224] = `IFUPATH806.swl.thr0_state;
thread_status[3225] = `IFUPATH806.swl.thr1_state;
thread_status[3226] = `IFUPATH806.swl.thr2_state;
thread_status[3227] = `IFUPATH806.swl.thr3_state;
thread_status[3228] = `IFUPATH807.swl.thr0_state;
thread_status[3229] = `IFUPATH807.swl.thr1_state;
thread_status[3230] = `IFUPATH807.swl.thr2_state;
thread_status[3231] = `IFUPATH807.swl.thr3_state;
thread_status[3232] = `IFUPATH808.swl.thr0_state;
thread_status[3233] = `IFUPATH808.swl.thr1_state;
thread_status[3234] = `IFUPATH808.swl.thr2_state;
thread_status[3235] = `IFUPATH808.swl.thr3_state;
thread_status[3236] = `IFUPATH809.swl.thr0_state;
thread_status[3237] = `IFUPATH809.swl.thr1_state;
thread_status[3238] = `IFUPATH809.swl.thr2_state;
thread_status[3239] = `IFUPATH809.swl.thr3_state;
thread_status[3240] = `IFUPATH810.swl.thr0_state;
thread_status[3241] = `IFUPATH810.swl.thr1_state;
thread_status[3242] = `IFUPATH810.swl.thr2_state;
thread_status[3243] = `IFUPATH810.swl.thr3_state;
thread_status[3244] = `IFUPATH811.swl.thr0_state;
thread_status[3245] = `IFUPATH811.swl.thr1_state;
thread_status[3246] = `IFUPATH811.swl.thr2_state;
thread_status[3247] = `IFUPATH811.swl.thr3_state;
thread_status[3248] = `IFUPATH812.swl.thr0_state;
thread_status[3249] = `IFUPATH812.swl.thr1_state;
thread_status[3250] = `IFUPATH812.swl.thr2_state;
thread_status[3251] = `IFUPATH812.swl.thr3_state;
thread_status[3252] = `IFUPATH813.swl.thr0_state;
thread_status[3253] = `IFUPATH813.swl.thr1_state;
thread_status[3254] = `IFUPATH813.swl.thr2_state;
thread_status[3255] = `IFUPATH813.swl.thr3_state;
thread_status[3256] = `IFUPATH814.swl.thr0_state;
thread_status[3257] = `IFUPATH814.swl.thr1_state;
thread_status[3258] = `IFUPATH814.swl.thr2_state;
thread_status[3259] = `IFUPATH814.swl.thr3_state;
thread_status[3260] = `IFUPATH815.swl.thr0_state;
thread_status[3261] = `IFUPATH815.swl.thr1_state;
thread_status[3262] = `IFUPATH815.swl.thr2_state;
thread_status[3263] = `IFUPATH815.swl.thr3_state;
thread_status[3264] = `IFUPATH816.swl.thr0_state;
thread_status[3265] = `IFUPATH816.swl.thr1_state;
thread_status[3266] = `IFUPATH816.swl.thr2_state;
thread_status[3267] = `IFUPATH816.swl.thr3_state;
thread_status[3268] = `IFUPATH817.swl.thr0_state;
thread_status[3269] = `IFUPATH817.swl.thr1_state;
thread_status[3270] = `IFUPATH817.swl.thr2_state;
thread_status[3271] = `IFUPATH817.swl.thr3_state;
thread_status[3272] = `IFUPATH818.swl.thr0_state;
thread_status[3273] = `IFUPATH818.swl.thr1_state;
thread_status[3274] = `IFUPATH818.swl.thr2_state;
thread_status[3275] = `IFUPATH818.swl.thr3_state;
thread_status[3276] = `IFUPATH819.swl.thr0_state;
thread_status[3277] = `IFUPATH819.swl.thr1_state;
thread_status[3278] = `IFUPATH819.swl.thr2_state;
thread_status[3279] = `IFUPATH819.swl.thr3_state;
thread_status[3280] = `IFUPATH820.swl.thr0_state;
thread_status[3281] = `IFUPATH820.swl.thr1_state;
thread_status[3282] = `IFUPATH820.swl.thr2_state;
thread_status[3283] = `IFUPATH820.swl.thr3_state;
thread_status[3284] = `IFUPATH821.swl.thr0_state;
thread_status[3285] = `IFUPATH821.swl.thr1_state;
thread_status[3286] = `IFUPATH821.swl.thr2_state;
thread_status[3287] = `IFUPATH821.swl.thr3_state;
thread_status[3288] = `IFUPATH822.swl.thr0_state;
thread_status[3289] = `IFUPATH822.swl.thr1_state;
thread_status[3290] = `IFUPATH822.swl.thr2_state;
thread_status[3291] = `IFUPATH822.swl.thr3_state;
thread_status[3292] = `IFUPATH823.swl.thr0_state;
thread_status[3293] = `IFUPATH823.swl.thr1_state;
thread_status[3294] = `IFUPATH823.swl.thr2_state;
thread_status[3295] = `IFUPATH823.swl.thr3_state;
thread_status[3296] = `IFUPATH824.swl.thr0_state;
thread_status[3297] = `IFUPATH824.swl.thr1_state;
thread_status[3298] = `IFUPATH824.swl.thr2_state;
thread_status[3299] = `IFUPATH824.swl.thr3_state;
thread_status[3300] = `IFUPATH825.swl.thr0_state;
thread_status[3301] = `IFUPATH825.swl.thr1_state;
thread_status[3302] = `IFUPATH825.swl.thr2_state;
thread_status[3303] = `IFUPATH825.swl.thr3_state;
thread_status[3304] = `IFUPATH826.swl.thr0_state;
thread_status[3305] = `IFUPATH826.swl.thr1_state;
thread_status[3306] = `IFUPATH826.swl.thr2_state;
thread_status[3307] = `IFUPATH826.swl.thr3_state;
thread_status[3308] = `IFUPATH827.swl.thr0_state;
thread_status[3309] = `IFUPATH827.swl.thr1_state;
thread_status[3310] = `IFUPATH827.swl.thr2_state;
thread_status[3311] = `IFUPATH827.swl.thr3_state;
thread_status[3312] = `IFUPATH828.swl.thr0_state;
thread_status[3313] = `IFUPATH828.swl.thr1_state;
thread_status[3314] = `IFUPATH828.swl.thr2_state;
thread_status[3315] = `IFUPATH828.swl.thr3_state;
thread_status[3316] = `IFUPATH829.swl.thr0_state;
thread_status[3317] = `IFUPATH829.swl.thr1_state;
thread_status[3318] = `IFUPATH829.swl.thr2_state;
thread_status[3319] = `IFUPATH829.swl.thr3_state;
thread_status[3320] = `IFUPATH830.swl.thr0_state;
thread_status[3321] = `IFUPATH830.swl.thr1_state;
thread_status[3322] = `IFUPATH830.swl.thr2_state;
thread_status[3323] = `IFUPATH830.swl.thr3_state;
thread_status[3324] = `IFUPATH831.swl.thr0_state;
thread_status[3325] = `IFUPATH831.swl.thr1_state;
thread_status[3326] = `IFUPATH831.swl.thr2_state;
thread_status[3327] = `IFUPATH831.swl.thr3_state;
thread_status[3328] = `IFUPATH832.swl.thr0_state;
thread_status[3329] = `IFUPATH832.swl.thr1_state;
thread_status[3330] = `IFUPATH832.swl.thr2_state;
thread_status[3331] = `IFUPATH832.swl.thr3_state;
thread_status[3332] = `IFUPATH833.swl.thr0_state;
thread_status[3333] = `IFUPATH833.swl.thr1_state;
thread_status[3334] = `IFUPATH833.swl.thr2_state;
thread_status[3335] = `IFUPATH833.swl.thr3_state;
thread_status[3336] = `IFUPATH834.swl.thr0_state;
thread_status[3337] = `IFUPATH834.swl.thr1_state;
thread_status[3338] = `IFUPATH834.swl.thr2_state;
thread_status[3339] = `IFUPATH834.swl.thr3_state;
thread_status[3340] = `IFUPATH835.swl.thr0_state;
thread_status[3341] = `IFUPATH835.swl.thr1_state;
thread_status[3342] = `IFUPATH835.swl.thr2_state;
thread_status[3343] = `IFUPATH835.swl.thr3_state;
thread_status[3344] = `IFUPATH836.swl.thr0_state;
thread_status[3345] = `IFUPATH836.swl.thr1_state;
thread_status[3346] = `IFUPATH836.swl.thr2_state;
thread_status[3347] = `IFUPATH836.swl.thr3_state;
thread_status[3348] = `IFUPATH837.swl.thr0_state;
thread_status[3349] = `IFUPATH837.swl.thr1_state;
thread_status[3350] = `IFUPATH837.swl.thr2_state;
thread_status[3351] = `IFUPATH837.swl.thr3_state;
thread_status[3352] = `IFUPATH838.swl.thr0_state;
thread_status[3353] = `IFUPATH838.swl.thr1_state;
thread_status[3354] = `IFUPATH838.swl.thr2_state;
thread_status[3355] = `IFUPATH838.swl.thr3_state;
thread_status[3356] = `IFUPATH839.swl.thr0_state;
thread_status[3357] = `IFUPATH839.swl.thr1_state;
thread_status[3358] = `IFUPATH839.swl.thr2_state;
thread_status[3359] = `IFUPATH839.swl.thr3_state;
thread_status[3360] = `IFUPATH840.swl.thr0_state;
thread_status[3361] = `IFUPATH840.swl.thr1_state;
thread_status[3362] = `IFUPATH840.swl.thr2_state;
thread_status[3363] = `IFUPATH840.swl.thr3_state;
thread_status[3364] = `IFUPATH841.swl.thr0_state;
thread_status[3365] = `IFUPATH841.swl.thr1_state;
thread_status[3366] = `IFUPATH841.swl.thr2_state;
thread_status[3367] = `IFUPATH841.swl.thr3_state;
thread_status[3368] = `IFUPATH842.swl.thr0_state;
thread_status[3369] = `IFUPATH842.swl.thr1_state;
thread_status[3370] = `IFUPATH842.swl.thr2_state;
thread_status[3371] = `IFUPATH842.swl.thr3_state;
thread_status[3372] = `IFUPATH843.swl.thr0_state;
thread_status[3373] = `IFUPATH843.swl.thr1_state;
thread_status[3374] = `IFUPATH843.swl.thr2_state;
thread_status[3375] = `IFUPATH843.swl.thr3_state;
thread_status[3376] = `IFUPATH844.swl.thr0_state;
thread_status[3377] = `IFUPATH844.swl.thr1_state;
thread_status[3378] = `IFUPATH844.swl.thr2_state;
thread_status[3379] = `IFUPATH844.swl.thr3_state;
thread_status[3380] = `IFUPATH845.swl.thr0_state;
thread_status[3381] = `IFUPATH845.swl.thr1_state;
thread_status[3382] = `IFUPATH845.swl.thr2_state;
thread_status[3383] = `IFUPATH845.swl.thr3_state;
thread_status[3384] = `IFUPATH846.swl.thr0_state;
thread_status[3385] = `IFUPATH846.swl.thr1_state;
thread_status[3386] = `IFUPATH846.swl.thr2_state;
thread_status[3387] = `IFUPATH846.swl.thr3_state;
thread_status[3388] = `IFUPATH847.swl.thr0_state;
thread_status[3389] = `IFUPATH847.swl.thr1_state;
thread_status[3390] = `IFUPATH847.swl.thr2_state;
thread_status[3391] = `IFUPATH847.swl.thr3_state;
thread_status[3392] = `IFUPATH848.swl.thr0_state;
thread_status[3393] = `IFUPATH848.swl.thr1_state;
thread_status[3394] = `IFUPATH848.swl.thr2_state;
thread_status[3395] = `IFUPATH848.swl.thr3_state;
thread_status[3396] = `IFUPATH849.swl.thr0_state;
thread_status[3397] = `IFUPATH849.swl.thr1_state;
thread_status[3398] = `IFUPATH849.swl.thr2_state;
thread_status[3399] = `IFUPATH849.swl.thr3_state;
thread_status[3400] = `IFUPATH850.swl.thr0_state;
thread_status[3401] = `IFUPATH850.swl.thr1_state;
thread_status[3402] = `IFUPATH850.swl.thr2_state;
thread_status[3403] = `IFUPATH850.swl.thr3_state;
thread_status[3404] = `IFUPATH851.swl.thr0_state;
thread_status[3405] = `IFUPATH851.swl.thr1_state;
thread_status[3406] = `IFUPATH851.swl.thr2_state;
thread_status[3407] = `IFUPATH851.swl.thr3_state;
thread_status[3408] = `IFUPATH852.swl.thr0_state;
thread_status[3409] = `IFUPATH852.swl.thr1_state;
thread_status[3410] = `IFUPATH852.swl.thr2_state;
thread_status[3411] = `IFUPATH852.swl.thr3_state;
thread_status[3412] = `IFUPATH853.swl.thr0_state;
thread_status[3413] = `IFUPATH853.swl.thr1_state;
thread_status[3414] = `IFUPATH853.swl.thr2_state;
thread_status[3415] = `IFUPATH853.swl.thr3_state;
thread_status[3416] = `IFUPATH854.swl.thr0_state;
thread_status[3417] = `IFUPATH854.swl.thr1_state;
thread_status[3418] = `IFUPATH854.swl.thr2_state;
thread_status[3419] = `IFUPATH854.swl.thr3_state;
thread_status[3420] = `IFUPATH855.swl.thr0_state;
thread_status[3421] = `IFUPATH855.swl.thr1_state;
thread_status[3422] = `IFUPATH855.swl.thr2_state;
thread_status[3423] = `IFUPATH855.swl.thr3_state;
thread_status[3424] = `IFUPATH856.swl.thr0_state;
thread_status[3425] = `IFUPATH856.swl.thr1_state;
thread_status[3426] = `IFUPATH856.swl.thr2_state;
thread_status[3427] = `IFUPATH856.swl.thr3_state;
thread_status[3428] = `IFUPATH857.swl.thr0_state;
thread_status[3429] = `IFUPATH857.swl.thr1_state;
thread_status[3430] = `IFUPATH857.swl.thr2_state;
thread_status[3431] = `IFUPATH857.swl.thr3_state;
thread_status[3432] = `IFUPATH858.swl.thr0_state;
thread_status[3433] = `IFUPATH858.swl.thr1_state;
thread_status[3434] = `IFUPATH858.swl.thr2_state;
thread_status[3435] = `IFUPATH858.swl.thr3_state;
thread_status[3436] = `IFUPATH859.swl.thr0_state;
thread_status[3437] = `IFUPATH859.swl.thr1_state;
thread_status[3438] = `IFUPATH859.swl.thr2_state;
thread_status[3439] = `IFUPATH859.swl.thr3_state;
thread_status[3440] = `IFUPATH860.swl.thr0_state;
thread_status[3441] = `IFUPATH860.swl.thr1_state;
thread_status[3442] = `IFUPATH860.swl.thr2_state;
thread_status[3443] = `IFUPATH860.swl.thr3_state;
thread_status[3444] = `IFUPATH861.swl.thr0_state;
thread_status[3445] = `IFUPATH861.swl.thr1_state;
thread_status[3446] = `IFUPATH861.swl.thr2_state;
thread_status[3447] = `IFUPATH861.swl.thr3_state;
thread_status[3448] = `IFUPATH862.swl.thr0_state;
thread_status[3449] = `IFUPATH862.swl.thr1_state;
thread_status[3450] = `IFUPATH862.swl.thr2_state;
thread_status[3451] = `IFUPATH862.swl.thr3_state;
thread_status[3452] = `IFUPATH863.swl.thr0_state;
thread_status[3453] = `IFUPATH863.swl.thr1_state;
thread_status[3454] = `IFUPATH863.swl.thr2_state;
thread_status[3455] = `IFUPATH863.swl.thr3_state;
thread_status[3456] = `IFUPATH864.swl.thr0_state;
thread_status[3457] = `IFUPATH864.swl.thr1_state;
thread_status[3458] = `IFUPATH864.swl.thr2_state;
thread_status[3459] = `IFUPATH864.swl.thr3_state;
thread_status[3460] = `IFUPATH865.swl.thr0_state;
thread_status[3461] = `IFUPATH865.swl.thr1_state;
thread_status[3462] = `IFUPATH865.swl.thr2_state;
thread_status[3463] = `IFUPATH865.swl.thr3_state;
thread_status[3464] = `IFUPATH866.swl.thr0_state;
thread_status[3465] = `IFUPATH866.swl.thr1_state;
thread_status[3466] = `IFUPATH866.swl.thr2_state;
thread_status[3467] = `IFUPATH866.swl.thr3_state;
thread_status[3468] = `IFUPATH867.swl.thr0_state;
thread_status[3469] = `IFUPATH867.swl.thr1_state;
thread_status[3470] = `IFUPATH867.swl.thr2_state;
thread_status[3471] = `IFUPATH867.swl.thr3_state;
thread_status[3472] = `IFUPATH868.swl.thr0_state;
thread_status[3473] = `IFUPATH868.swl.thr1_state;
thread_status[3474] = `IFUPATH868.swl.thr2_state;
thread_status[3475] = `IFUPATH868.swl.thr3_state;
thread_status[3476] = `IFUPATH869.swl.thr0_state;
thread_status[3477] = `IFUPATH869.swl.thr1_state;
thread_status[3478] = `IFUPATH869.swl.thr2_state;
thread_status[3479] = `IFUPATH869.swl.thr3_state;
thread_status[3480] = `IFUPATH870.swl.thr0_state;
thread_status[3481] = `IFUPATH870.swl.thr1_state;
thread_status[3482] = `IFUPATH870.swl.thr2_state;
thread_status[3483] = `IFUPATH870.swl.thr3_state;
thread_status[3484] = `IFUPATH871.swl.thr0_state;
thread_status[3485] = `IFUPATH871.swl.thr1_state;
thread_status[3486] = `IFUPATH871.swl.thr2_state;
thread_status[3487] = `IFUPATH871.swl.thr3_state;
thread_status[3488] = `IFUPATH872.swl.thr0_state;
thread_status[3489] = `IFUPATH872.swl.thr1_state;
thread_status[3490] = `IFUPATH872.swl.thr2_state;
thread_status[3491] = `IFUPATH872.swl.thr3_state;
thread_status[3492] = `IFUPATH873.swl.thr0_state;
thread_status[3493] = `IFUPATH873.swl.thr1_state;
thread_status[3494] = `IFUPATH873.swl.thr2_state;
thread_status[3495] = `IFUPATH873.swl.thr3_state;
thread_status[3496] = `IFUPATH874.swl.thr0_state;
thread_status[3497] = `IFUPATH874.swl.thr1_state;
thread_status[3498] = `IFUPATH874.swl.thr2_state;
thread_status[3499] = `IFUPATH874.swl.thr3_state;
thread_status[3500] = `IFUPATH875.swl.thr0_state;
thread_status[3501] = `IFUPATH875.swl.thr1_state;
thread_status[3502] = `IFUPATH875.swl.thr2_state;
thread_status[3503] = `IFUPATH875.swl.thr3_state;
thread_status[3504] = `IFUPATH876.swl.thr0_state;
thread_status[3505] = `IFUPATH876.swl.thr1_state;
thread_status[3506] = `IFUPATH876.swl.thr2_state;
thread_status[3507] = `IFUPATH876.swl.thr3_state;
thread_status[3508] = `IFUPATH877.swl.thr0_state;
thread_status[3509] = `IFUPATH877.swl.thr1_state;
thread_status[3510] = `IFUPATH877.swl.thr2_state;
thread_status[3511] = `IFUPATH877.swl.thr3_state;
thread_status[3512] = `IFUPATH878.swl.thr0_state;
thread_status[3513] = `IFUPATH878.swl.thr1_state;
thread_status[3514] = `IFUPATH878.swl.thr2_state;
thread_status[3515] = `IFUPATH878.swl.thr3_state;
thread_status[3516] = `IFUPATH879.swl.thr0_state;
thread_status[3517] = `IFUPATH879.swl.thr1_state;
thread_status[3518] = `IFUPATH879.swl.thr2_state;
thread_status[3519] = `IFUPATH879.swl.thr3_state;
thread_status[3520] = `IFUPATH880.swl.thr0_state;
thread_status[3521] = `IFUPATH880.swl.thr1_state;
thread_status[3522] = `IFUPATH880.swl.thr2_state;
thread_status[3523] = `IFUPATH880.swl.thr3_state;
thread_status[3524] = `IFUPATH881.swl.thr0_state;
thread_status[3525] = `IFUPATH881.swl.thr1_state;
thread_status[3526] = `IFUPATH881.swl.thr2_state;
thread_status[3527] = `IFUPATH881.swl.thr3_state;
thread_status[3528] = `IFUPATH882.swl.thr0_state;
thread_status[3529] = `IFUPATH882.swl.thr1_state;
thread_status[3530] = `IFUPATH882.swl.thr2_state;
thread_status[3531] = `IFUPATH882.swl.thr3_state;
thread_status[3532] = `IFUPATH883.swl.thr0_state;
thread_status[3533] = `IFUPATH883.swl.thr1_state;
thread_status[3534] = `IFUPATH883.swl.thr2_state;
thread_status[3535] = `IFUPATH883.swl.thr3_state;
thread_status[3536] = `IFUPATH884.swl.thr0_state;
thread_status[3537] = `IFUPATH884.swl.thr1_state;
thread_status[3538] = `IFUPATH884.swl.thr2_state;
thread_status[3539] = `IFUPATH884.swl.thr3_state;
thread_status[3540] = `IFUPATH885.swl.thr0_state;
thread_status[3541] = `IFUPATH885.swl.thr1_state;
thread_status[3542] = `IFUPATH885.swl.thr2_state;
thread_status[3543] = `IFUPATH885.swl.thr3_state;
thread_status[3544] = `IFUPATH886.swl.thr0_state;
thread_status[3545] = `IFUPATH886.swl.thr1_state;
thread_status[3546] = `IFUPATH886.swl.thr2_state;
thread_status[3547] = `IFUPATH886.swl.thr3_state;
thread_status[3548] = `IFUPATH887.swl.thr0_state;
thread_status[3549] = `IFUPATH887.swl.thr1_state;
thread_status[3550] = `IFUPATH887.swl.thr2_state;
thread_status[3551] = `IFUPATH887.swl.thr3_state;
thread_status[3552] = `IFUPATH888.swl.thr0_state;
thread_status[3553] = `IFUPATH888.swl.thr1_state;
thread_status[3554] = `IFUPATH888.swl.thr2_state;
thread_status[3555] = `IFUPATH888.swl.thr3_state;
thread_status[3556] = `IFUPATH889.swl.thr0_state;
thread_status[3557] = `IFUPATH889.swl.thr1_state;
thread_status[3558] = `IFUPATH889.swl.thr2_state;
thread_status[3559] = `IFUPATH889.swl.thr3_state;
thread_status[3560] = `IFUPATH890.swl.thr0_state;
thread_status[3561] = `IFUPATH890.swl.thr1_state;
thread_status[3562] = `IFUPATH890.swl.thr2_state;
thread_status[3563] = `IFUPATH890.swl.thr3_state;
thread_status[3564] = `IFUPATH891.swl.thr0_state;
thread_status[3565] = `IFUPATH891.swl.thr1_state;
thread_status[3566] = `IFUPATH891.swl.thr2_state;
thread_status[3567] = `IFUPATH891.swl.thr3_state;
thread_status[3568] = `IFUPATH892.swl.thr0_state;
thread_status[3569] = `IFUPATH892.swl.thr1_state;
thread_status[3570] = `IFUPATH892.swl.thr2_state;
thread_status[3571] = `IFUPATH892.swl.thr3_state;
thread_status[3572] = `IFUPATH893.swl.thr0_state;
thread_status[3573] = `IFUPATH893.swl.thr1_state;
thread_status[3574] = `IFUPATH893.swl.thr2_state;
thread_status[3575] = `IFUPATH893.swl.thr3_state;
thread_status[3576] = `IFUPATH894.swl.thr0_state;
thread_status[3577] = `IFUPATH894.swl.thr1_state;
thread_status[3578] = `IFUPATH894.swl.thr2_state;
thread_status[3579] = `IFUPATH894.swl.thr3_state;
thread_status[3580] = `IFUPATH895.swl.thr0_state;
thread_status[3581] = `IFUPATH895.swl.thr1_state;
thread_status[3582] = `IFUPATH895.swl.thr2_state;
thread_status[3583] = `IFUPATH895.swl.thr3_state;
thread_status[3584] = `IFUPATH896.swl.thr0_state;
thread_status[3585] = `IFUPATH896.swl.thr1_state;
thread_status[3586] = `IFUPATH896.swl.thr2_state;
thread_status[3587] = `IFUPATH896.swl.thr3_state;
thread_status[3588] = `IFUPATH897.swl.thr0_state;
thread_status[3589] = `IFUPATH897.swl.thr1_state;
thread_status[3590] = `IFUPATH897.swl.thr2_state;
thread_status[3591] = `IFUPATH897.swl.thr3_state;
thread_status[3592] = `IFUPATH898.swl.thr0_state;
thread_status[3593] = `IFUPATH898.swl.thr1_state;
thread_status[3594] = `IFUPATH898.swl.thr2_state;
thread_status[3595] = `IFUPATH898.swl.thr3_state;
thread_status[3596] = `IFUPATH899.swl.thr0_state;
thread_status[3597] = `IFUPATH899.swl.thr1_state;
thread_status[3598] = `IFUPATH899.swl.thr2_state;
thread_status[3599] = `IFUPATH899.swl.thr3_state;
thread_status[3600] = `IFUPATH900.swl.thr0_state;
thread_status[3601] = `IFUPATH900.swl.thr1_state;
thread_status[3602] = `IFUPATH900.swl.thr2_state;
thread_status[3603] = `IFUPATH900.swl.thr3_state;
thread_status[3604] = `IFUPATH901.swl.thr0_state;
thread_status[3605] = `IFUPATH901.swl.thr1_state;
thread_status[3606] = `IFUPATH901.swl.thr2_state;
thread_status[3607] = `IFUPATH901.swl.thr3_state;
thread_status[3608] = `IFUPATH902.swl.thr0_state;
thread_status[3609] = `IFUPATH902.swl.thr1_state;
thread_status[3610] = `IFUPATH902.swl.thr2_state;
thread_status[3611] = `IFUPATH902.swl.thr3_state;
thread_status[3612] = `IFUPATH903.swl.thr0_state;
thread_status[3613] = `IFUPATH903.swl.thr1_state;
thread_status[3614] = `IFUPATH903.swl.thr2_state;
thread_status[3615] = `IFUPATH903.swl.thr3_state;
thread_status[3616] = `IFUPATH904.swl.thr0_state;
thread_status[3617] = `IFUPATH904.swl.thr1_state;
thread_status[3618] = `IFUPATH904.swl.thr2_state;
thread_status[3619] = `IFUPATH904.swl.thr3_state;
thread_status[3620] = `IFUPATH905.swl.thr0_state;
thread_status[3621] = `IFUPATH905.swl.thr1_state;
thread_status[3622] = `IFUPATH905.swl.thr2_state;
thread_status[3623] = `IFUPATH905.swl.thr3_state;
thread_status[3624] = `IFUPATH906.swl.thr0_state;
thread_status[3625] = `IFUPATH906.swl.thr1_state;
thread_status[3626] = `IFUPATH906.swl.thr2_state;
thread_status[3627] = `IFUPATH906.swl.thr3_state;
thread_status[3628] = `IFUPATH907.swl.thr0_state;
thread_status[3629] = `IFUPATH907.swl.thr1_state;
thread_status[3630] = `IFUPATH907.swl.thr2_state;
thread_status[3631] = `IFUPATH907.swl.thr3_state;
thread_status[3632] = `IFUPATH908.swl.thr0_state;
thread_status[3633] = `IFUPATH908.swl.thr1_state;
thread_status[3634] = `IFUPATH908.swl.thr2_state;
thread_status[3635] = `IFUPATH908.swl.thr3_state;
thread_status[3636] = `IFUPATH909.swl.thr0_state;
thread_status[3637] = `IFUPATH909.swl.thr1_state;
thread_status[3638] = `IFUPATH909.swl.thr2_state;
thread_status[3639] = `IFUPATH909.swl.thr3_state;
thread_status[3640] = `IFUPATH910.swl.thr0_state;
thread_status[3641] = `IFUPATH910.swl.thr1_state;
thread_status[3642] = `IFUPATH910.swl.thr2_state;
thread_status[3643] = `IFUPATH910.swl.thr3_state;
thread_status[3644] = `IFUPATH911.swl.thr0_state;
thread_status[3645] = `IFUPATH911.swl.thr1_state;
thread_status[3646] = `IFUPATH911.swl.thr2_state;
thread_status[3647] = `IFUPATH911.swl.thr3_state;
thread_status[3648] = `IFUPATH912.swl.thr0_state;
thread_status[3649] = `IFUPATH912.swl.thr1_state;
thread_status[3650] = `IFUPATH912.swl.thr2_state;
thread_status[3651] = `IFUPATH912.swl.thr3_state;
thread_status[3652] = `IFUPATH913.swl.thr0_state;
thread_status[3653] = `IFUPATH913.swl.thr1_state;
thread_status[3654] = `IFUPATH913.swl.thr2_state;
thread_status[3655] = `IFUPATH913.swl.thr3_state;
thread_status[3656] = `IFUPATH914.swl.thr0_state;
thread_status[3657] = `IFUPATH914.swl.thr1_state;
thread_status[3658] = `IFUPATH914.swl.thr2_state;
thread_status[3659] = `IFUPATH914.swl.thr3_state;
thread_status[3660] = `IFUPATH915.swl.thr0_state;
thread_status[3661] = `IFUPATH915.swl.thr1_state;
thread_status[3662] = `IFUPATH915.swl.thr2_state;
thread_status[3663] = `IFUPATH915.swl.thr3_state;
thread_status[3664] = `IFUPATH916.swl.thr0_state;
thread_status[3665] = `IFUPATH916.swl.thr1_state;
thread_status[3666] = `IFUPATH916.swl.thr2_state;
thread_status[3667] = `IFUPATH916.swl.thr3_state;
thread_status[3668] = `IFUPATH917.swl.thr0_state;
thread_status[3669] = `IFUPATH917.swl.thr1_state;
thread_status[3670] = `IFUPATH917.swl.thr2_state;
thread_status[3671] = `IFUPATH917.swl.thr3_state;
thread_status[3672] = `IFUPATH918.swl.thr0_state;
thread_status[3673] = `IFUPATH918.swl.thr1_state;
thread_status[3674] = `IFUPATH918.swl.thr2_state;
thread_status[3675] = `IFUPATH918.swl.thr3_state;
thread_status[3676] = `IFUPATH919.swl.thr0_state;
thread_status[3677] = `IFUPATH919.swl.thr1_state;
thread_status[3678] = `IFUPATH919.swl.thr2_state;
thread_status[3679] = `IFUPATH919.swl.thr3_state;
thread_status[3680] = `IFUPATH920.swl.thr0_state;
thread_status[3681] = `IFUPATH920.swl.thr1_state;
thread_status[3682] = `IFUPATH920.swl.thr2_state;
thread_status[3683] = `IFUPATH920.swl.thr3_state;
thread_status[3684] = `IFUPATH921.swl.thr0_state;
thread_status[3685] = `IFUPATH921.swl.thr1_state;
thread_status[3686] = `IFUPATH921.swl.thr2_state;
thread_status[3687] = `IFUPATH921.swl.thr3_state;
thread_status[3688] = `IFUPATH922.swl.thr0_state;
thread_status[3689] = `IFUPATH922.swl.thr1_state;
thread_status[3690] = `IFUPATH922.swl.thr2_state;
thread_status[3691] = `IFUPATH922.swl.thr3_state;
thread_status[3692] = `IFUPATH923.swl.thr0_state;
thread_status[3693] = `IFUPATH923.swl.thr1_state;
thread_status[3694] = `IFUPATH923.swl.thr2_state;
thread_status[3695] = `IFUPATH923.swl.thr3_state;
thread_status[3696] = `IFUPATH924.swl.thr0_state;
thread_status[3697] = `IFUPATH924.swl.thr1_state;
thread_status[3698] = `IFUPATH924.swl.thr2_state;
thread_status[3699] = `IFUPATH924.swl.thr3_state;
thread_status[3700] = `IFUPATH925.swl.thr0_state;
thread_status[3701] = `IFUPATH925.swl.thr1_state;
thread_status[3702] = `IFUPATH925.swl.thr2_state;
thread_status[3703] = `IFUPATH925.swl.thr3_state;
thread_status[3704] = `IFUPATH926.swl.thr0_state;
thread_status[3705] = `IFUPATH926.swl.thr1_state;
thread_status[3706] = `IFUPATH926.swl.thr2_state;
thread_status[3707] = `IFUPATH926.swl.thr3_state;
thread_status[3708] = `IFUPATH927.swl.thr0_state;
thread_status[3709] = `IFUPATH927.swl.thr1_state;
thread_status[3710] = `IFUPATH927.swl.thr2_state;
thread_status[3711] = `IFUPATH927.swl.thr3_state;
thread_status[3712] = `IFUPATH928.swl.thr0_state;
thread_status[3713] = `IFUPATH928.swl.thr1_state;
thread_status[3714] = `IFUPATH928.swl.thr2_state;
thread_status[3715] = `IFUPATH928.swl.thr3_state;
thread_status[3716] = `IFUPATH929.swl.thr0_state;
thread_status[3717] = `IFUPATH929.swl.thr1_state;
thread_status[3718] = `IFUPATH929.swl.thr2_state;
thread_status[3719] = `IFUPATH929.swl.thr3_state;
thread_status[3720] = `IFUPATH930.swl.thr0_state;
thread_status[3721] = `IFUPATH930.swl.thr1_state;
thread_status[3722] = `IFUPATH930.swl.thr2_state;
thread_status[3723] = `IFUPATH930.swl.thr3_state;
thread_status[3724] = `IFUPATH931.swl.thr0_state;
thread_status[3725] = `IFUPATH931.swl.thr1_state;
thread_status[3726] = `IFUPATH931.swl.thr2_state;
thread_status[3727] = `IFUPATH931.swl.thr3_state;
thread_status[3728] = `IFUPATH932.swl.thr0_state;
thread_status[3729] = `IFUPATH932.swl.thr1_state;
thread_status[3730] = `IFUPATH932.swl.thr2_state;
thread_status[3731] = `IFUPATH932.swl.thr3_state;
thread_status[3732] = `IFUPATH933.swl.thr0_state;
thread_status[3733] = `IFUPATH933.swl.thr1_state;
thread_status[3734] = `IFUPATH933.swl.thr2_state;
thread_status[3735] = `IFUPATH933.swl.thr3_state;
thread_status[3736] = `IFUPATH934.swl.thr0_state;
thread_status[3737] = `IFUPATH934.swl.thr1_state;
thread_status[3738] = `IFUPATH934.swl.thr2_state;
thread_status[3739] = `IFUPATH934.swl.thr3_state;
thread_status[3740] = `IFUPATH935.swl.thr0_state;
thread_status[3741] = `IFUPATH935.swl.thr1_state;
thread_status[3742] = `IFUPATH935.swl.thr2_state;
thread_status[3743] = `IFUPATH935.swl.thr3_state;
thread_status[3744] = `IFUPATH936.swl.thr0_state;
thread_status[3745] = `IFUPATH936.swl.thr1_state;
thread_status[3746] = `IFUPATH936.swl.thr2_state;
thread_status[3747] = `IFUPATH936.swl.thr3_state;
thread_status[3748] = `IFUPATH937.swl.thr0_state;
thread_status[3749] = `IFUPATH937.swl.thr1_state;
thread_status[3750] = `IFUPATH937.swl.thr2_state;
thread_status[3751] = `IFUPATH937.swl.thr3_state;
thread_status[3752] = `IFUPATH938.swl.thr0_state;
thread_status[3753] = `IFUPATH938.swl.thr1_state;
thread_status[3754] = `IFUPATH938.swl.thr2_state;
thread_status[3755] = `IFUPATH938.swl.thr3_state;
thread_status[3756] = `IFUPATH939.swl.thr0_state;
thread_status[3757] = `IFUPATH939.swl.thr1_state;
thread_status[3758] = `IFUPATH939.swl.thr2_state;
thread_status[3759] = `IFUPATH939.swl.thr3_state;
thread_status[3760] = `IFUPATH940.swl.thr0_state;
thread_status[3761] = `IFUPATH940.swl.thr1_state;
thread_status[3762] = `IFUPATH940.swl.thr2_state;
thread_status[3763] = `IFUPATH940.swl.thr3_state;
thread_status[3764] = `IFUPATH941.swl.thr0_state;
thread_status[3765] = `IFUPATH941.swl.thr1_state;
thread_status[3766] = `IFUPATH941.swl.thr2_state;
thread_status[3767] = `IFUPATH941.swl.thr3_state;
thread_status[3768] = `IFUPATH942.swl.thr0_state;
thread_status[3769] = `IFUPATH942.swl.thr1_state;
thread_status[3770] = `IFUPATH942.swl.thr2_state;
thread_status[3771] = `IFUPATH942.swl.thr3_state;
thread_status[3772] = `IFUPATH943.swl.thr0_state;
thread_status[3773] = `IFUPATH943.swl.thr1_state;
thread_status[3774] = `IFUPATH943.swl.thr2_state;
thread_status[3775] = `IFUPATH943.swl.thr3_state;
thread_status[3776] = `IFUPATH944.swl.thr0_state;
thread_status[3777] = `IFUPATH944.swl.thr1_state;
thread_status[3778] = `IFUPATH944.swl.thr2_state;
thread_status[3779] = `IFUPATH944.swl.thr3_state;
thread_status[3780] = `IFUPATH945.swl.thr0_state;
thread_status[3781] = `IFUPATH945.swl.thr1_state;
thread_status[3782] = `IFUPATH945.swl.thr2_state;
thread_status[3783] = `IFUPATH945.swl.thr3_state;
thread_status[3784] = `IFUPATH946.swl.thr0_state;
thread_status[3785] = `IFUPATH946.swl.thr1_state;
thread_status[3786] = `IFUPATH946.swl.thr2_state;
thread_status[3787] = `IFUPATH946.swl.thr3_state;
thread_status[3788] = `IFUPATH947.swl.thr0_state;
thread_status[3789] = `IFUPATH947.swl.thr1_state;
thread_status[3790] = `IFUPATH947.swl.thr2_state;
thread_status[3791] = `IFUPATH947.swl.thr3_state;
thread_status[3792] = `IFUPATH948.swl.thr0_state;
thread_status[3793] = `IFUPATH948.swl.thr1_state;
thread_status[3794] = `IFUPATH948.swl.thr2_state;
thread_status[3795] = `IFUPATH948.swl.thr3_state;
thread_status[3796] = `IFUPATH949.swl.thr0_state;
thread_status[3797] = `IFUPATH949.swl.thr1_state;
thread_status[3798] = `IFUPATH949.swl.thr2_state;
thread_status[3799] = `IFUPATH949.swl.thr3_state;
thread_status[3800] = `IFUPATH950.swl.thr0_state;
thread_status[3801] = `IFUPATH950.swl.thr1_state;
thread_status[3802] = `IFUPATH950.swl.thr2_state;
thread_status[3803] = `IFUPATH950.swl.thr3_state;
thread_status[3804] = `IFUPATH951.swl.thr0_state;
thread_status[3805] = `IFUPATH951.swl.thr1_state;
thread_status[3806] = `IFUPATH951.swl.thr2_state;
thread_status[3807] = `IFUPATH951.swl.thr3_state;
thread_status[3808] = `IFUPATH952.swl.thr0_state;
thread_status[3809] = `IFUPATH952.swl.thr1_state;
thread_status[3810] = `IFUPATH952.swl.thr2_state;
thread_status[3811] = `IFUPATH952.swl.thr3_state;
thread_status[3812] = `IFUPATH953.swl.thr0_state;
thread_status[3813] = `IFUPATH953.swl.thr1_state;
thread_status[3814] = `IFUPATH953.swl.thr2_state;
thread_status[3815] = `IFUPATH953.swl.thr3_state;
thread_status[3816] = `IFUPATH954.swl.thr0_state;
thread_status[3817] = `IFUPATH954.swl.thr1_state;
thread_status[3818] = `IFUPATH954.swl.thr2_state;
thread_status[3819] = `IFUPATH954.swl.thr3_state;
thread_status[3820] = `IFUPATH955.swl.thr0_state;
thread_status[3821] = `IFUPATH955.swl.thr1_state;
thread_status[3822] = `IFUPATH955.swl.thr2_state;
thread_status[3823] = `IFUPATH955.swl.thr3_state;
thread_status[3824] = `IFUPATH956.swl.thr0_state;
thread_status[3825] = `IFUPATH956.swl.thr1_state;
thread_status[3826] = `IFUPATH956.swl.thr2_state;
thread_status[3827] = `IFUPATH956.swl.thr3_state;
thread_status[3828] = `IFUPATH957.swl.thr0_state;
thread_status[3829] = `IFUPATH957.swl.thr1_state;
thread_status[3830] = `IFUPATH957.swl.thr2_state;
thread_status[3831] = `IFUPATH957.swl.thr3_state;
thread_status[3832] = `IFUPATH958.swl.thr0_state;
thread_status[3833] = `IFUPATH958.swl.thr1_state;
thread_status[3834] = `IFUPATH958.swl.thr2_state;
thread_status[3835] = `IFUPATH958.swl.thr3_state;
thread_status[3836] = `IFUPATH959.swl.thr0_state;
thread_status[3837] = `IFUPATH959.swl.thr1_state;
thread_status[3838] = `IFUPATH959.swl.thr2_state;
thread_status[3839] = `IFUPATH959.swl.thr3_state;
thread_status[3840] = `IFUPATH960.swl.thr0_state;
thread_status[3841] = `IFUPATH960.swl.thr1_state;
thread_status[3842] = `IFUPATH960.swl.thr2_state;
thread_status[3843] = `IFUPATH960.swl.thr3_state;
thread_status[3844] = `IFUPATH961.swl.thr0_state;
thread_status[3845] = `IFUPATH961.swl.thr1_state;
thread_status[3846] = `IFUPATH961.swl.thr2_state;
thread_status[3847] = `IFUPATH961.swl.thr3_state;
thread_status[3848] = `IFUPATH962.swl.thr0_state;
thread_status[3849] = `IFUPATH962.swl.thr1_state;
thread_status[3850] = `IFUPATH962.swl.thr2_state;
thread_status[3851] = `IFUPATH962.swl.thr3_state;
thread_status[3852] = `IFUPATH963.swl.thr0_state;
thread_status[3853] = `IFUPATH963.swl.thr1_state;
thread_status[3854] = `IFUPATH963.swl.thr2_state;
thread_status[3855] = `IFUPATH963.swl.thr3_state;
thread_status[3856] = `IFUPATH964.swl.thr0_state;
thread_status[3857] = `IFUPATH964.swl.thr1_state;
thread_status[3858] = `IFUPATH964.swl.thr2_state;
thread_status[3859] = `IFUPATH964.swl.thr3_state;
thread_status[3860] = `IFUPATH965.swl.thr0_state;
thread_status[3861] = `IFUPATH965.swl.thr1_state;
thread_status[3862] = `IFUPATH965.swl.thr2_state;
thread_status[3863] = `IFUPATH965.swl.thr3_state;
thread_status[3864] = `IFUPATH966.swl.thr0_state;
thread_status[3865] = `IFUPATH966.swl.thr1_state;
thread_status[3866] = `IFUPATH966.swl.thr2_state;
thread_status[3867] = `IFUPATH966.swl.thr3_state;
thread_status[3868] = `IFUPATH967.swl.thr0_state;
thread_status[3869] = `IFUPATH967.swl.thr1_state;
thread_status[3870] = `IFUPATH967.swl.thr2_state;
thread_status[3871] = `IFUPATH967.swl.thr3_state;
thread_status[3872] = `IFUPATH968.swl.thr0_state;
thread_status[3873] = `IFUPATH968.swl.thr1_state;
thread_status[3874] = `IFUPATH968.swl.thr2_state;
thread_status[3875] = `IFUPATH968.swl.thr3_state;
thread_status[3876] = `IFUPATH969.swl.thr0_state;
thread_status[3877] = `IFUPATH969.swl.thr1_state;
thread_status[3878] = `IFUPATH969.swl.thr2_state;
thread_status[3879] = `IFUPATH969.swl.thr3_state;
thread_status[3880] = `IFUPATH970.swl.thr0_state;
thread_status[3881] = `IFUPATH970.swl.thr1_state;
thread_status[3882] = `IFUPATH970.swl.thr2_state;
thread_status[3883] = `IFUPATH970.swl.thr3_state;
thread_status[3884] = `IFUPATH971.swl.thr0_state;
thread_status[3885] = `IFUPATH971.swl.thr1_state;
thread_status[3886] = `IFUPATH971.swl.thr2_state;
thread_status[3887] = `IFUPATH971.swl.thr3_state;
thread_status[3888] = `IFUPATH972.swl.thr0_state;
thread_status[3889] = `IFUPATH972.swl.thr1_state;
thread_status[3890] = `IFUPATH972.swl.thr2_state;
thread_status[3891] = `IFUPATH972.swl.thr3_state;
thread_status[3892] = `IFUPATH973.swl.thr0_state;
thread_status[3893] = `IFUPATH973.swl.thr1_state;
thread_status[3894] = `IFUPATH973.swl.thr2_state;
thread_status[3895] = `IFUPATH973.swl.thr3_state;
thread_status[3896] = `IFUPATH974.swl.thr0_state;
thread_status[3897] = `IFUPATH974.swl.thr1_state;
thread_status[3898] = `IFUPATH974.swl.thr2_state;
thread_status[3899] = `IFUPATH974.swl.thr3_state;
thread_status[3900] = `IFUPATH975.swl.thr0_state;
thread_status[3901] = `IFUPATH975.swl.thr1_state;
thread_status[3902] = `IFUPATH975.swl.thr2_state;
thread_status[3903] = `IFUPATH975.swl.thr3_state;
thread_status[3904] = `IFUPATH976.swl.thr0_state;
thread_status[3905] = `IFUPATH976.swl.thr1_state;
thread_status[3906] = `IFUPATH976.swl.thr2_state;
thread_status[3907] = `IFUPATH976.swl.thr3_state;
thread_status[3908] = `IFUPATH977.swl.thr0_state;
thread_status[3909] = `IFUPATH977.swl.thr1_state;
thread_status[3910] = `IFUPATH977.swl.thr2_state;
thread_status[3911] = `IFUPATH977.swl.thr3_state;
thread_status[3912] = `IFUPATH978.swl.thr0_state;
thread_status[3913] = `IFUPATH978.swl.thr1_state;
thread_status[3914] = `IFUPATH978.swl.thr2_state;
thread_status[3915] = `IFUPATH978.swl.thr3_state;
thread_status[3916] = `IFUPATH979.swl.thr0_state;
thread_status[3917] = `IFUPATH979.swl.thr1_state;
thread_status[3918] = `IFUPATH979.swl.thr2_state;
thread_status[3919] = `IFUPATH979.swl.thr3_state;
thread_status[3920] = `IFUPATH980.swl.thr0_state;
thread_status[3921] = `IFUPATH980.swl.thr1_state;
thread_status[3922] = `IFUPATH980.swl.thr2_state;
thread_status[3923] = `IFUPATH980.swl.thr3_state;
thread_status[3924] = `IFUPATH981.swl.thr0_state;
thread_status[3925] = `IFUPATH981.swl.thr1_state;
thread_status[3926] = `IFUPATH981.swl.thr2_state;
thread_status[3927] = `IFUPATH981.swl.thr3_state;
thread_status[3928] = `IFUPATH982.swl.thr0_state;
thread_status[3929] = `IFUPATH982.swl.thr1_state;
thread_status[3930] = `IFUPATH982.swl.thr2_state;
thread_status[3931] = `IFUPATH982.swl.thr3_state;
thread_status[3932] = `IFUPATH983.swl.thr0_state;
thread_status[3933] = `IFUPATH983.swl.thr1_state;
thread_status[3934] = `IFUPATH983.swl.thr2_state;
thread_status[3935] = `IFUPATH983.swl.thr3_state;
thread_status[3936] = `IFUPATH984.swl.thr0_state;
thread_status[3937] = `IFUPATH984.swl.thr1_state;
thread_status[3938] = `IFUPATH984.swl.thr2_state;
thread_status[3939] = `IFUPATH984.swl.thr3_state;
thread_status[3940] = `IFUPATH985.swl.thr0_state;
thread_status[3941] = `IFUPATH985.swl.thr1_state;
thread_status[3942] = `IFUPATH985.swl.thr2_state;
thread_status[3943] = `IFUPATH985.swl.thr3_state;
thread_status[3944] = `IFUPATH986.swl.thr0_state;
thread_status[3945] = `IFUPATH986.swl.thr1_state;
thread_status[3946] = `IFUPATH986.swl.thr2_state;
thread_status[3947] = `IFUPATH986.swl.thr3_state;
thread_status[3948] = `IFUPATH987.swl.thr0_state;
thread_status[3949] = `IFUPATH987.swl.thr1_state;
thread_status[3950] = `IFUPATH987.swl.thr2_state;
thread_status[3951] = `IFUPATH987.swl.thr3_state;
thread_status[3952] = `IFUPATH988.swl.thr0_state;
thread_status[3953] = `IFUPATH988.swl.thr1_state;
thread_status[3954] = `IFUPATH988.swl.thr2_state;
thread_status[3955] = `IFUPATH988.swl.thr3_state;
thread_status[3956] = `IFUPATH989.swl.thr0_state;
thread_status[3957] = `IFUPATH989.swl.thr1_state;
thread_status[3958] = `IFUPATH989.swl.thr2_state;
thread_status[3959] = `IFUPATH989.swl.thr3_state;
thread_status[3960] = `IFUPATH990.swl.thr0_state;
thread_status[3961] = `IFUPATH990.swl.thr1_state;
thread_status[3962] = `IFUPATH990.swl.thr2_state;
thread_status[3963] = `IFUPATH990.swl.thr3_state;
thread_status[3964] = `IFUPATH991.swl.thr0_state;
thread_status[3965] = `IFUPATH991.swl.thr1_state;
thread_status[3966] = `IFUPATH991.swl.thr2_state;
thread_status[3967] = `IFUPATH991.swl.thr3_state;
thread_status[3968] = `IFUPATH992.swl.thr0_state;
thread_status[3969] = `IFUPATH992.swl.thr1_state;
thread_status[3970] = `IFUPATH992.swl.thr2_state;
thread_status[3971] = `IFUPATH992.swl.thr3_state;
thread_status[3972] = `IFUPATH993.swl.thr0_state;
thread_status[3973] = `IFUPATH993.swl.thr1_state;
thread_status[3974] = `IFUPATH993.swl.thr2_state;
thread_status[3975] = `IFUPATH993.swl.thr3_state;
thread_status[3976] = `IFUPATH994.swl.thr0_state;
thread_status[3977] = `IFUPATH994.swl.thr1_state;
thread_status[3978] = `IFUPATH994.swl.thr2_state;
thread_status[3979] = `IFUPATH994.swl.thr3_state;
thread_status[3980] = `IFUPATH995.swl.thr0_state;
thread_status[3981] = `IFUPATH995.swl.thr1_state;
thread_status[3982] = `IFUPATH995.swl.thr2_state;
thread_status[3983] = `IFUPATH995.swl.thr3_state;
thread_status[3984] = `IFUPATH996.swl.thr0_state;
thread_status[3985] = `IFUPATH996.swl.thr1_state;
thread_status[3986] = `IFUPATH996.swl.thr2_state;
thread_status[3987] = `IFUPATH996.swl.thr3_state;
thread_status[3988] = `IFUPATH997.swl.thr0_state;
thread_status[3989] = `IFUPATH997.swl.thr1_state;
thread_status[3990] = `IFUPATH997.swl.thr2_state;
thread_status[3991] = `IFUPATH997.swl.thr3_state;
thread_status[3992] = `IFUPATH998.swl.thr0_state;
thread_status[3993] = `IFUPATH998.swl.thr1_state;
thread_status[3994] = `IFUPATH998.swl.thr2_state;
thread_status[3995] = `IFUPATH998.swl.thr3_state;
thread_status[3996] = `IFUPATH999.swl.thr0_state;
thread_status[3997] = `IFUPATH999.swl.thr1_state;
thread_status[3998] = `IFUPATH999.swl.thr2_state;
thread_status[3999] = `IFUPATH999.swl.thr3_state;
thread_status[4000] = `IFUPATH1000.swl.thr0_state;
thread_status[4001] = `IFUPATH1000.swl.thr1_state;
thread_status[4002] = `IFUPATH1000.swl.thr2_state;
thread_status[4003] = `IFUPATH1000.swl.thr3_state;
thread_status[4004] = `IFUPATH1001.swl.thr0_state;
thread_status[4005] = `IFUPATH1001.swl.thr1_state;
thread_status[4006] = `IFUPATH1001.swl.thr2_state;
thread_status[4007] = `IFUPATH1001.swl.thr3_state;
thread_status[4008] = `IFUPATH1002.swl.thr0_state;
thread_status[4009] = `IFUPATH1002.swl.thr1_state;
thread_status[4010] = `IFUPATH1002.swl.thr2_state;
thread_status[4011] = `IFUPATH1002.swl.thr3_state;
thread_status[4012] = `IFUPATH1003.swl.thr0_state;
thread_status[4013] = `IFUPATH1003.swl.thr1_state;
thread_status[4014] = `IFUPATH1003.swl.thr2_state;
thread_status[4015] = `IFUPATH1003.swl.thr3_state;
thread_status[4016] = `IFUPATH1004.swl.thr0_state;
thread_status[4017] = `IFUPATH1004.swl.thr1_state;
thread_status[4018] = `IFUPATH1004.swl.thr2_state;
thread_status[4019] = `IFUPATH1004.swl.thr3_state;
thread_status[4020] = `IFUPATH1005.swl.thr0_state;
thread_status[4021] = `IFUPATH1005.swl.thr1_state;
thread_status[4022] = `IFUPATH1005.swl.thr2_state;
thread_status[4023] = `IFUPATH1005.swl.thr3_state;
thread_status[4024] = `IFUPATH1006.swl.thr0_state;
thread_status[4025] = `IFUPATH1006.swl.thr1_state;
thread_status[4026] = `IFUPATH1006.swl.thr2_state;
thread_status[4027] = `IFUPATH1006.swl.thr3_state;
thread_status[4028] = `IFUPATH1007.swl.thr0_state;
thread_status[4029] = `IFUPATH1007.swl.thr1_state;
thread_status[4030] = `IFUPATH1007.swl.thr2_state;
thread_status[4031] = `IFUPATH1007.swl.thr3_state;
thread_status[4032] = `IFUPATH1008.swl.thr0_state;
thread_status[4033] = `IFUPATH1008.swl.thr1_state;
thread_status[4034] = `IFUPATH1008.swl.thr2_state;
thread_status[4035] = `IFUPATH1008.swl.thr3_state;
thread_status[4036] = `IFUPATH1009.swl.thr0_state;
thread_status[4037] = `IFUPATH1009.swl.thr1_state;
thread_status[4038] = `IFUPATH1009.swl.thr2_state;
thread_status[4039] = `IFUPATH1009.swl.thr3_state;
thread_status[4040] = `IFUPATH1010.swl.thr0_state;
thread_status[4041] = `IFUPATH1010.swl.thr1_state;
thread_status[4042] = `IFUPATH1010.swl.thr2_state;
thread_status[4043] = `IFUPATH1010.swl.thr3_state;
thread_status[4044] = `IFUPATH1011.swl.thr0_state;
thread_status[4045] = `IFUPATH1011.swl.thr1_state;
thread_status[4046] = `IFUPATH1011.swl.thr2_state;
thread_status[4047] = `IFUPATH1011.swl.thr3_state;
thread_status[4048] = `IFUPATH1012.swl.thr0_state;
thread_status[4049] = `IFUPATH1012.swl.thr1_state;
thread_status[4050] = `IFUPATH1012.swl.thr2_state;
thread_status[4051] = `IFUPATH1012.swl.thr3_state;
thread_status[4052] = `IFUPATH1013.swl.thr0_state;
thread_status[4053] = `IFUPATH1013.swl.thr1_state;
thread_status[4054] = `IFUPATH1013.swl.thr2_state;
thread_status[4055] = `IFUPATH1013.swl.thr3_state;
thread_status[4056] = `IFUPATH1014.swl.thr0_state;
thread_status[4057] = `IFUPATH1014.swl.thr1_state;
thread_status[4058] = `IFUPATH1014.swl.thr2_state;
thread_status[4059] = `IFUPATH1014.swl.thr3_state;
thread_status[4060] = `IFUPATH1015.swl.thr0_state;
thread_status[4061] = `IFUPATH1015.swl.thr1_state;
thread_status[4062] = `IFUPATH1015.swl.thr2_state;
thread_status[4063] = `IFUPATH1015.swl.thr3_state;
thread_status[4064] = `IFUPATH1016.swl.thr0_state;
thread_status[4065] = `IFUPATH1016.swl.thr1_state;
thread_status[4066] = `IFUPATH1016.swl.thr2_state;
thread_status[4067] = `IFUPATH1016.swl.thr3_state;
thread_status[4068] = `IFUPATH1017.swl.thr0_state;
thread_status[4069] = `IFUPATH1017.swl.thr1_state;
thread_status[4070] = `IFUPATH1017.swl.thr2_state;
thread_status[4071] = `IFUPATH1017.swl.thr3_state;
thread_status[4072] = `IFUPATH1018.swl.thr0_state;
thread_status[4073] = `IFUPATH1018.swl.thr1_state;
thread_status[4074] = `IFUPATH1018.swl.thr2_state;
thread_status[4075] = `IFUPATH1018.swl.thr3_state;
thread_status[4076] = `IFUPATH1019.swl.thr0_state;
thread_status[4077] = `IFUPATH1019.swl.thr1_state;
thread_status[4078] = `IFUPATH1019.swl.thr2_state;
thread_status[4079] = `IFUPATH1019.swl.thr3_state;
thread_status[4080] = `IFUPATH1020.swl.thr0_state;
thread_status[4081] = `IFUPATH1020.swl.thr1_state;
thread_status[4082] = `IFUPATH1020.swl.thr2_state;
thread_status[4083] = `IFUPATH1020.swl.thr3_state;
thread_status[4084] = `IFUPATH1021.swl.thr0_state;
thread_status[4085] = `IFUPATH1021.swl.thr1_state;
thread_status[4086] = `IFUPATH1021.swl.thr2_state;
thread_status[4087] = `IFUPATH1021.swl.thr3_state;
thread_status[4088] = `IFUPATH1022.swl.thr0_state;
thread_status[4089] = `IFUPATH1022.swl.thr1_state;
thread_status[4090] = `IFUPATH1022.swl.thr2_state;
thread_status[4091] = `IFUPATH1022.swl.thr3_state;
thread_status[4092] = `IFUPATH1023.swl.thr0_state;
thread_status[4093] = `IFUPATH1023.swl.thr1_state;
thread_status[4094] = `IFUPATH1023.swl.thr2_state;
thread_status[4095] = `IFUPATH1023.swl.thr3_state;

    end
endtask // get_thread_status
`endif


            assign spc0_thread_id = 2'b00;
            assign spc0_rtl_pc = spc0_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(0*4)]   <= 1'b0;
                  active_thread[(0*4)+1] <= 1'b0;
                  active_thread[(0*4)+2] <= 1'b0;
                  active_thread[(0*4)+3] <= 1'b0;
                  spc0_inst_done         <= 0;
                  spc0_phy_pc_w          <= 0;
                end else begin
                  active_thread[(0*4)]   <= 1'b1;
                  active_thread[(0*4)+1] <= 1'b1;
                  active_thread[(0*4)+2] <= 1'b1;
                  active_thread[(0*4)+3] <= 1'b1;
                  spc0_inst_done         <= `ARIANE_CORE0.piton_pc_vld;
                  spc0_phy_pc_w          <= `ARIANE_CORE0.piton_pc;
                end
            end
    

            assign spc1_thread_id = 2'b00;
            assign spc1_rtl_pc = spc1_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(1*4)]   <= 1'b0;
                  active_thread[(1*4)+1] <= 1'b0;
                  active_thread[(1*4)+2] <= 1'b0;
                  active_thread[(1*4)+3] <= 1'b0;
                  spc1_inst_done         <= 0;
                  spc1_phy_pc_w          <= 0;
                end else begin
                  active_thread[(1*4)]   <= 1'b1;
                  active_thread[(1*4)+1] <= 1'b1;
                  active_thread[(1*4)+2] <= 1'b1;
                  active_thread[(1*4)+3] <= 1'b1;
                  spc1_inst_done         <= `ARIANE_CORE1.piton_pc_vld;
                  spc1_phy_pc_w          <= `ARIANE_CORE1.piton_pc;
                end
            end
    

            assign spc2_thread_id = 2'b00;
            assign spc2_rtl_pc = spc2_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(2*4)]   <= 1'b0;
                  active_thread[(2*4)+1] <= 1'b0;
                  active_thread[(2*4)+2] <= 1'b0;
                  active_thread[(2*4)+3] <= 1'b0;
                  spc2_inst_done         <= 0;
                  spc2_phy_pc_w          <= 0;
                end else begin
                  active_thread[(2*4)]   <= 1'b1;
                  active_thread[(2*4)+1] <= 1'b1;
                  active_thread[(2*4)+2] <= 1'b1;
                  active_thread[(2*4)+3] <= 1'b1;
                  spc2_inst_done         <= `ARIANE_CORE2.piton_pc_vld;
                  spc2_phy_pc_w          <= `ARIANE_CORE2.piton_pc;
                end
            end
    

            assign spc3_thread_id = 2'b00;
            assign spc3_rtl_pc = spc3_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(3*4)]   <= 1'b0;
                  active_thread[(3*4)+1] <= 1'b0;
                  active_thread[(3*4)+2] <= 1'b0;
                  active_thread[(3*4)+3] <= 1'b0;
                  spc3_inst_done         <= 0;
                  spc3_phy_pc_w          <= 0;
                end else begin
                  active_thread[(3*4)]   <= 1'b1;
                  active_thread[(3*4)+1] <= 1'b1;
                  active_thread[(3*4)+2] <= 1'b1;
                  active_thread[(3*4)+3] <= 1'b1;
                  spc3_inst_done         <= `ARIANE_CORE3.piton_pc_vld;
                  spc3_phy_pc_w          <= `ARIANE_CORE3.piton_pc;
                end
            end
    

            assign spc4_thread_id = 2'b00;
            assign spc4_rtl_pc = spc4_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(4*4)]   <= 1'b0;
                  active_thread[(4*4)+1] <= 1'b0;
                  active_thread[(4*4)+2] <= 1'b0;
                  active_thread[(4*4)+3] <= 1'b0;
                  spc4_inst_done         <= 0;
                  spc4_phy_pc_w          <= 0;
                end else begin
                  active_thread[(4*4)]   <= 1'b1;
                  active_thread[(4*4)+1] <= 1'b1;
                  active_thread[(4*4)+2] <= 1'b1;
                  active_thread[(4*4)+3] <= 1'b1;
                  spc4_inst_done         <= `ARIANE_CORE4.piton_pc_vld;
                  spc4_phy_pc_w          <= `ARIANE_CORE4.piton_pc;
                end
            end
    

            assign spc5_thread_id = 2'b00;
            assign spc5_rtl_pc = spc5_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(5*4)]   <= 1'b0;
                  active_thread[(5*4)+1] <= 1'b0;
                  active_thread[(5*4)+2] <= 1'b0;
                  active_thread[(5*4)+3] <= 1'b0;
                  spc5_inst_done         <= 0;
                  spc5_phy_pc_w          <= 0;
                end else begin
                  active_thread[(5*4)]   <= 1'b1;
                  active_thread[(5*4)+1] <= 1'b1;
                  active_thread[(5*4)+2] <= 1'b1;
                  active_thread[(5*4)+3] <= 1'b1;
                  spc5_inst_done         <= `ARIANE_CORE5.piton_pc_vld;
                  spc5_phy_pc_w          <= `ARIANE_CORE5.piton_pc;
                end
            end
    

            assign spc6_thread_id = 2'b00;
            assign spc6_rtl_pc = spc6_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(6*4)]   <= 1'b0;
                  active_thread[(6*4)+1] <= 1'b0;
                  active_thread[(6*4)+2] <= 1'b0;
                  active_thread[(6*4)+3] <= 1'b0;
                  spc6_inst_done         <= 0;
                  spc6_phy_pc_w          <= 0;
                end else begin
                  active_thread[(6*4)]   <= 1'b1;
                  active_thread[(6*4)+1] <= 1'b1;
                  active_thread[(6*4)+2] <= 1'b1;
                  active_thread[(6*4)+3] <= 1'b1;
                  spc6_inst_done         <= `ARIANE_CORE6.piton_pc_vld;
                  spc6_phy_pc_w          <= `ARIANE_CORE6.piton_pc;
                end
            end
    

            assign spc7_thread_id = 2'b00;
            assign spc7_rtl_pc = spc7_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(7*4)]   <= 1'b0;
                  active_thread[(7*4)+1] <= 1'b0;
                  active_thread[(7*4)+2] <= 1'b0;
                  active_thread[(7*4)+3] <= 1'b0;
                  spc7_inst_done         <= 0;
                  spc7_phy_pc_w          <= 0;
                end else begin
                  active_thread[(7*4)]   <= 1'b1;
                  active_thread[(7*4)+1] <= 1'b1;
                  active_thread[(7*4)+2] <= 1'b1;
                  active_thread[(7*4)+3] <= 1'b1;
                  spc7_inst_done         <= `ARIANE_CORE7.piton_pc_vld;
                  spc7_phy_pc_w          <= `ARIANE_CORE7.piton_pc;
                end
            end
    

            assign spc8_thread_id = 2'b00;
            assign spc8_rtl_pc = spc8_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(8*4)]   <= 1'b0;
                  active_thread[(8*4)+1] <= 1'b0;
                  active_thread[(8*4)+2] <= 1'b0;
                  active_thread[(8*4)+3] <= 1'b0;
                  spc8_inst_done         <= 0;
                  spc8_phy_pc_w          <= 0;
                end else begin
                  active_thread[(8*4)]   <= 1'b1;
                  active_thread[(8*4)+1] <= 1'b1;
                  active_thread[(8*4)+2] <= 1'b1;
                  active_thread[(8*4)+3] <= 1'b1;
                  spc8_inst_done         <= `ARIANE_CORE8.piton_pc_vld;
                  spc8_phy_pc_w          <= `ARIANE_CORE8.piton_pc;
                end
            end
    

            assign spc9_thread_id = 2'b00;
            assign spc9_rtl_pc = spc9_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(9*4)]   <= 1'b0;
                  active_thread[(9*4)+1] <= 1'b0;
                  active_thread[(9*4)+2] <= 1'b0;
                  active_thread[(9*4)+3] <= 1'b0;
                  spc9_inst_done         <= 0;
                  spc9_phy_pc_w          <= 0;
                end else begin
                  active_thread[(9*4)]   <= 1'b1;
                  active_thread[(9*4)+1] <= 1'b1;
                  active_thread[(9*4)+2] <= 1'b1;
                  active_thread[(9*4)+3] <= 1'b1;
                  spc9_inst_done         <= `ARIANE_CORE9.piton_pc_vld;
                  spc9_phy_pc_w          <= `ARIANE_CORE9.piton_pc;
                end
            end
    

            assign spc10_thread_id = 2'b00;
            assign spc10_rtl_pc = spc10_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(10*4)]   <= 1'b0;
                  active_thread[(10*4)+1] <= 1'b0;
                  active_thread[(10*4)+2] <= 1'b0;
                  active_thread[(10*4)+3] <= 1'b0;
                  spc10_inst_done         <= 0;
                  spc10_phy_pc_w          <= 0;
                end else begin
                  active_thread[(10*4)]   <= 1'b1;
                  active_thread[(10*4)+1] <= 1'b1;
                  active_thread[(10*4)+2] <= 1'b1;
                  active_thread[(10*4)+3] <= 1'b1;
                  spc10_inst_done         <= `ARIANE_CORE10.piton_pc_vld;
                  spc10_phy_pc_w          <= `ARIANE_CORE10.piton_pc;
                end
            end
    

            assign spc11_thread_id = 2'b00;
            assign spc11_rtl_pc = spc11_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(11*4)]   <= 1'b0;
                  active_thread[(11*4)+1] <= 1'b0;
                  active_thread[(11*4)+2] <= 1'b0;
                  active_thread[(11*4)+3] <= 1'b0;
                  spc11_inst_done         <= 0;
                  spc11_phy_pc_w          <= 0;
                end else begin
                  active_thread[(11*4)]   <= 1'b1;
                  active_thread[(11*4)+1] <= 1'b1;
                  active_thread[(11*4)+2] <= 1'b1;
                  active_thread[(11*4)+3] <= 1'b1;
                  spc11_inst_done         <= `ARIANE_CORE11.piton_pc_vld;
                  spc11_phy_pc_w          <= `ARIANE_CORE11.piton_pc;
                end
            end
    

            assign spc12_thread_id = 2'b00;
            assign spc12_rtl_pc = spc12_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(12*4)]   <= 1'b0;
                  active_thread[(12*4)+1] <= 1'b0;
                  active_thread[(12*4)+2] <= 1'b0;
                  active_thread[(12*4)+3] <= 1'b0;
                  spc12_inst_done         <= 0;
                  spc12_phy_pc_w          <= 0;
                end else begin
                  active_thread[(12*4)]   <= 1'b1;
                  active_thread[(12*4)+1] <= 1'b1;
                  active_thread[(12*4)+2] <= 1'b1;
                  active_thread[(12*4)+3] <= 1'b1;
                  spc12_inst_done         <= `ARIANE_CORE12.piton_pc_vld;
                  spc12_phy_pc_w          <= `ARIANE_CORE12.piton_pc;
                end
            end
    

            assign spc13_thread_id = 2'b00;
            assign spc13_rtl_pc = spc13_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(13*4)]   <= 1'b0;
                  active_thread[(13*4)+1] <= 1'b0;
                  active_thread[(13*4)+2] <= 1'b0;
                  active_thread[(13*4)+3] <= 1'b0;
                  spc13_inst_done         <= 0;
                  spc13_phy_pc_w          <= 0;
                end else begin
                  active_thread[(13*4)]   <= 1'b1;
                  active_thread[(13*4)+1] <= 1'b1;
                  active_thread[(13*4)+2] <= 1'b1;
                  active_thread[(13*4)+3] <= 1'b1;
                  spc13_inst_done         <= `ARIANE_CORE13.piton_pc_vld;
                  spc13_phy_pc_w          <= `ARIANE_CORE13.piton_pc;
                end
            end
    

            assign spc14_thread_id = 2'b00;
            assign spc14_rtl_pc = spc14_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(14*4)]   <= 1'b0;
                  active_thread[(14*4)+1] <= 1'b0;
                  active_thread[(14*4)+2] <= 1'b0;
                  active_thread[(14*4)+3] <= 1'b0;
                  spc14_inst_done         <= 0;
                  spc14_phy_pc_w          <= 0;
                end else begin
                  active_thread[(14*4)]   <= 1'b1;
                  active_thread[(14*4)+1] <= 1'b1;
                  active_thread[(14*4)+2] <= 1'b1;
                  active_thread[(14*4)+3] <= 1'b1;
                  spc14_inst_done         <= `ARIANE_CORE14.piton_pc_vld;
                  spc14_phy_pc_w          <= `ARIANE_CORE14.piton_pc;
                end
            end
    

            assign spc15_thread_id = 2'b00;
            assign spc15_rtl_pc = spc15_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(15*4)]   <= 1'b0;
                  active_thread[(15*4)+1] <= 1'b0;
                  active_thread[(15*4)+2] <= 1'b0;
                  active_thread[(15*4)+3] <= 1'b0;
                  spc15_inst_done         <= 0;
                  spc15_phy_pc_w          <= 0;
                end else begin
                  active_thread[(15*4)]   <= 1'b1;
                  active_thread[(15*4)+1] <= 1'b1;
                  active_thread[(15*4)+2] <= 1'b1;
                  active_thread[(15*4)+3] <= 1'b1;
                  spc15_inst_done         <= `ARIANE_CORE15.piton_pc_vld;
                  spc15_phy_pc_w          <= `ARIANE_CORE15.piton_pc;
                end
            end
    

            assign spc16_thread_id = 2'b00;
            assign spc16_rtl_pc = spc16_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(16*4)]   <= 1'b0;
                  active_thread[(16*4)+1] <= 1'b0;
                  active_thread[(16*4)+2] <= 1'b0;
                  active_thread[(16*4)+3] <= 1'b0;
                  spc16_inst_done         <= 0;
                  spc16_phy_pc_w          <= 0;
                end else begin
                  active_thread[(16*4)]   <= 1'b1;
                  active_thread[(16*4)+1] <= 1'b1;
                  active_thread[(16*4)+2] <= 1'b1;
                  active_thread[(16*4)+3] <= 1'b1;
                  spc16_inst_done         <= `ARIANE_CORE16.piton_pc_vld;
                  spc16_phy_pc_w          <= `ARIANE_CORE16.piton_pc;
                end
            end
    

            assign spc17_thread_id = 2'b00;
            assign spc17_rtl_pc = spc17_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(17*4)]   <= 1'b0;
                  active_thread[(17*4)+1] <= 1'b0;
                  active_thread[(17*4)+2] <= 1'b0;
                  active_thread[(17*4)+3] <= 1'b0;
                  spc17_inst_done         <= 0;
                  spc17_phy_pc_w          <= 0;
                end else begin
                  active_thread[(17*4)]   <= 1'b1;
                  active_thread[(17*4)+1] <= 1'b1;
                  active_thread[(17*4)+2] <= 1'b1;
                  active_thread[(17*4)+3] <= 1'b1;
                  spc17_inst_done         <= `ARIANE_CORE17.piton_pc_vld;
                  spc17_phy_pc_w          <= `ARIANE_CORE17.piton_pc;
                end
            end
    

            assign spc18_thread_id = 2'b00;
            assign spc18_rtl_pc = spc18_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(18*4)]   <= 1'b0;
                  active_thread[(18*4)+1] <= 1'b0;
                  active_thread[(18*4)+2] <= 1'b0;
                  active_thread[(18*4)+3] <= 1'b0;
                  spc18_inst_done         <= 0;
                  spc18_phy_pc_w          <= 0;
                end else begin
                  active_thread[(18*4)]   <= 1'b1;
                  active_thread[(18*4)+1] <= 1'b1;
                  active_thread[(18*4)+2] <= 1'b1;
                  active_thread[(18*4)+3] <= 1'b1;
                  spc18_inst_done         <= `ARIANE_CORE18.piton_pc_vld;
                  spc18_phy_pc_w          <= `ARIANE_CORE18.piton_pc;
                end
            end
    

            assign spc19_thread_id = 2'b00;
            assign spc19_rtl_pc = spc19_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(19*4)]   <= 1'b0;
                  active_thread[(19*4)+1] <= 1'b0;
                  active_thread[(19*4)+2] <= 1'b0;
                  active_thread[(19*4)+3] <= 1'b0;
                  spc19_inst_done         <= 0;
                  spc19_phy_pc_w          <= 0;
                end else begin
                  active_thread[(19*4)]   <= 1'b1;
                  active_thread[(19*4)+1] <= 1'b1;
                  active_thread[(19*4)+2] <= 1'b1;
                  active_thread[(19*4)+3] <= 1'b1;
                  spc19_inst_done         <= `ARIANE_CORE19.piton_pc_vld;
                  spc19_phy_pc_w          <= `ARIANE_CORE19.piton_pc;
                end
            end
    

            assign spc20_thread_id = 2'b00;
            assign spc20_rtl_pc = spc20_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(20*4)]   <= 1'b0;
                  active_thread[(20*4)+1] <= 1'b0;
                  active_thread[(20*4)+2] <= 1'b0;
                  active_thread[(20*4)+3] <= 1'b0;
                  spc20_inst_done         <= 0;
                  spc20_phy_pc_w          <= 0;
                end else begin
                  active_thread[(20*4)]   <= 1'b1;
                  active_thread[(20*4)+1] <= 1'b1;
                  active_thread[(20*4)+2] <= 1'b1;
                  active_thread[(20*4)+3] <= 1'b1;
                  spc20_inst_done         <= `ARIANE_CORE20.piton_pc_vld;
                  spc20_phy_pc_w          <= `ARIANE_CORE20.piton_pc;
                end
            end
    

            assign spc21_thread_id = 2'b00;
            assign spc21_rtl_pc = spc21_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(21*4)]   <= 1'b0;
                  active_thread[(21*4)+1] <= 1'b0;
                  active_thread[(21*4)+2] <= 1'b0;
                  active_thread[(21*4)+3] <= 1'b0;
                  spc21_inst_done         <= 0;
                  spc21_phy_pc_w          <= 0;
                end else begin
                  active_thread[(21*4)]   <= 1'b1;
                  active_thread[(21*4)+1] <= 1'b1;
                  active_thread[(21*4)+2] <= 1'b1;
                  active_thread[(21*4)+3] <= 1'b1;
                  spc21_inst_done         <= `ARIANE_CORE21.piton_pc_vld;
                  spc21_phy_pc_w          <= `ARIANE_CORE21.piton_pc;
                end
            end
    

            assign spc22_thread_id = 2'b00;
            assign spc22_rtl_pc = spc22_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(22*4)]   <= 1'b0;
                  active_thread[(22*4)+1] <= 1'b0;
                  active_thread[(22*4)+2] <= 1'b0;
                  active_thread[(22*4)+3] <= 1'b0;
                  spc22_inst_done         <= 0;
                  spc22_phy_pc_w          <= 0;
                end else begin
                  active_thread[(22*4)]   <= 1'b1;
                  active_thread[(22*4)+1] <= 1'b1;
                  active_thread[(22*4)+2] <= 1'b1;
                  active_thread[(22*4)+3] <= 1'b1;
                  spc22_inst_done         <= `ARIANE_CORE22.piton_pc_vld;
                  spc22_phy_pc_w          <= `ARIANE_CORE22.piton_pc;
                end
            end
    

            assign spc23_thread_id = 2'b00;
            assign spc23_rtl_pc = spc23_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(23*4)]   <= 1'b0;
                  active_thread[(23*4)+1] <= 1'b0;
                  active_thread[(23*4)+2] <= 1'b0;
                  active_thread[(23*4)+3] <= 1'b0;
                  spc23_inst_done         <= 0;
                  spc23_phy_pc_w          <= 0;
                end else begin
                  active_thread[(23*4)]   <= 1'b1;
                  active_thread[(23*4)+1] <= 1'b1;
                  active_thread[(23*4)+2] <= 1'b1;
                  active_thread[(23*4)+3] <= 1'b1;
                  spc23_inst_done         <= `ARIANE_CORE23.piton_pc_vld;
                  spc23_phy_pc_w          <= `ARIANE_CORE23.piton_pc;
                end
            end
    

            assign spc24_thread_id = 2'b00;
            assign spc24_rtl_pc = spc24_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(24*4)]   <= 1'b0;
                  active_thread[(24*4)+1] <= 1'b0;
                  active_thread[(24*4)+2] <= 1'b0;
                  active_thread[(24*4)+3] <= 1'b0;
                  spc24_inst_done         <= 0;
                  spc24_phy_pc_w          <= 0;
                end else begin
                  active_thread[(24*4)]   <= 1'b1;
                  active_thread[(24*4)+1] <= 1'b1;
                  active_thread[(24*4)+2] <= 1'b1;
                  active_thread[(24*4)+3] <= 1'b1;
                  spc24_inst_done         <= `ARIANE_CORE24.piton_pc_vld;
                  spc24_phy_pc_w          <= `ARIANE_CORE24.piton_pc;
                end
            end
    

            assign spc25_thread_id = 2'b00;
            assign spc25_rtl_pc = spc25_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(25*4)]   <= 1'b0;
                  active_thread[(25*4)+1] <= 1'b0;
                  active_thread[(25*4)+2] <= 1'b0;
                  active_thread[(25*4)+3] <= 1'b0;
                  spc25_inst_done         <= 0;
                  spc25_phy_pc_w          <= 0;
                end else begin
                  active_thread[(25*4)]   <= 1'b1;
                  active_thread[(25*4)+1] <= 1'b1;
                  active_thread[(25*4)+2] <= 1'b1;
                  active_thread[(25*4)+3] <= 1'b1;
                  spc25_inst_done         <= `ARIANE_CORE25.piton_pc_vld;
                  spc25_phy_pc_w          <= `ARIANE_CORE25.piton_pc;
                end
            end
    

            assign spc26_thread_id = 2'b00;
            assign spc26_rtl_pc = spc26_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(26*4)]   <= 1'b0;
                  active_thread[(26*4)+1] <= 1'b0;
                  active_thread[(26*4)+2] <= 1'b0;
                  active_thread[(26*4)+3] <= 1'b0;
                  spc26_inst_done         <= 0;
                  spc26_phy_pc_w          <= 0;
                end else begin
                  active_thread[(26*4)]   <= 1'b1;
                  active_thread[(26*4)+1] <= 1'b1;
                  active_thread[(26*4)+2] <= 1'b1;
                  active_thread[(26*4)+3] <= 1'b1;
                  spc26_inst_done         <= `ARIANE_CORE26.piton_pc_vld;
                  spc26_phy_pc_w          <= `ARIANE_CORE26.piton_pc;
                end
            end
    

            assign spc27_thread_id = 2'b00;
            assign spc27_rtl_pc = spc27_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(27*4)]   <= 1'b0;
                  active_thread[(27*4)+1] <= 1'b0;
                  active_thread[(27*4)+2] <= 1'b0;
                  active_thread[(27*4)+3] <= 1'b0;
                  spc27_inst_done         <= 0;
                  spc27_phy_pc_w          <= 0;
                end else begin
                  active_thread[(27*4)]   <= 1'b1;
                  active_thread[(27*4)+1] <= 1'b1;
                  active_thread[(27*4)+2] <= 1'b1;
                  active_thread[(27*4)+3] <= 1'b1;
                  spc27_inst_done         <= `ARIANE_CORE27.piton_pc_vld;
                  spc27_phy_pc_w          <= `ARIANE_CORE27.piton_pc;
                end
            end
    

            assign spc28_thread_id = 2'b00;
            assign spc28_rtl_pc = spc28_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(28*4)]   <= 1'b0;
                  active_thread[(28*4)+1] <= 1'b0;
                  active_thread[(28*4)+2] <= 1'b0;
                  active_thread[(28*4)+3] <= 1'b0;
                  spc28_inst_done         <= 0;
                  spc28_phy_pc_w          <= 0;
                end else begin
                  active_thread[(28*4)]   <= 1'b1;
                  active_thread[(28*4)+1] <= 1'b1;
                  active_thread[(28*4)+2] <= 1'b1;
                  active_thread[(28*4)+3] <= 1'b1;
                  spc28_inst_done         <= `ARIANE_CORE28.piton_pc_vld;
                  spc28_phy_pc_w          <= `ARIANE_CORE28.piton_pc;
                end
            end
    

            assign spc29_thread_id = 2'b00;
            assign spc29_rtl_pc = spc29_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(29*4)]   <= 1'b0;
                  active_thread[(29*4)+1] <= 1'b0;
                  active_thread[(29*4)+2] <= 1'b0;
                  active_thread[(29*4)+3] <= 1'b0;
                  spc29_inst_done         <= 0;
                  spc29_phy_pc_w          <= 0;
                end else begin
                  active_thread[(29*4)]   <= 1'b1;
                  active_thread[(29*4)+1] <= 1'b1;
                  active_thread[(29*4)+2] <= 1'b1;
                  active_thread[(29*4)+3] <= 1'b1;
                  spc29_inst_done         <= `ARIANE_CORE29.piton_pc_vld;
                  spc29_phy_pc_w          <= `ARIANE_CORE29.piton_pc;
                end
            end
    

            assign spc30_thread_id = 2'b00;
            assign spc30_rtl_pc = spc30_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(30*4)]   <= 1'b0;
                  active_thread[(30*4)+1] <= 1'b0;
                  active_thread[(30*4)+2] <= 1'b0;
                  active_thread[(30*4)+3] <= 1'b0;
                  spc30_inst_done         <= 0;
                  spc30_phy_pc_w          <= 0;
                end else begin
                  active_thread[(30*4)]   <= 1'b1;
                  active_thread[(30*4)+1] <= 1'b1;
                  active_thread[(30*4)+2] <= 1'b1;
                  active_thread[(30*4)+3] <= 1'b1;
                  spc30_inst_done         <= `ARIANE_CORE30.piton_pc_vld;
                  spc30_phy_pc_w          <= `ARIANE_CORE30.piton_pc;
                end
            end
    

            assign spc31_thread_id = 2'b00;
            assign spc31_rtl_pc = spc31_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(31*4)]   <= 1'b0;
                  active_thread[(31*4)+1] <= 1'b0;
                  active_thread[(31*4)+2] <= 1'b0;
                  active_thread[(31*4)+3] <= 1'b0;
                  spc31_inst_done         <= 0;
                  spc31_phy_pc_w          <= 0;
                end else begin
                  active_thread[(31*4)]   <= 1'b1;
                  active_thread[(31*4)+1] <= 1'b1;
                  active_thread[(31*4)+2] <= 1'b1;
                  active_thread[(31*4)+3] <= 1'b1;
                  spc31_inst_done         <= `ARIANE_CORE31.piton_pc_vld;
                  spc31_phy_pc_w          <= `ARIANE_CORE31.piton_pc;
                end
            end
    

            assign spc32_thread_id = 2'b00;
            assign spc32_rtl_pc = spc32_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(32*4)]   <= 1'b0;
                  active_thread[(32*4)+1] <= 1'b0;
                  active_thread[(32*4)+2] <= 1'b0;
                  active_thread[(32*4)+3] <= 1'b0;
                  spc32_inst_done         <= 0;
                  spc32_phy_pc_w          <= 0;
                end else begin
                  active_thread[(32*4)]   <= 1'b1;
                  active_thread[(32*4)+1] <= 1'b1;
                  active_thread[(32*4)+2] <= 1'b1;
                  active_thread[(32*4)+3] <= 1'b1;
                  spc32_inst_done         <= `ARIANE_CORE32.piton_pc_vld;
                  spc32_phy_pc_w          <= `ARIANE_CORE32.piton_pc;
                end
            end
    

            assign spc33_thread_id = 2'b00;
            assign spc33_rtl_pc = spc33_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(33*4)]   <= 1'b0;
                  active_thread[(33*4)+1] <= 1'b0;
                  active_thread[(33*4)+2] <= 1'b0;
                  active_thread[(33*4)+3] <= 1'b0;
                  spc33_inst_done         <= 0;
                  spc33_phy_pc_w          <= 0;
                end else begin
                  active_thread[(33*4)]   <= 1'b1;
                  active_thread[(33*4)+1] <= 1'b1;
                  active_thread[(33*4)+2] <= 1'b1;
                  active_thread[(33*4)+3] <= 1'b1;
                  spc33_inst_done         <= `ARIANE_CORE33.piton_pc_vld;
                  spc33_phy_pc_w          <= `ARIANE_CORE33.piton_pc;
                end
            end
    

            assign spc34_thread_id = 2'b00;
            assign spc34_rtl_pc = spc34_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(34*4)]   <= 1'b0;
                  active_thread[(34*4)+1] <= 1'b0;
                  active_thread[(34*4)+2] <= 1'b0;
                  active_thread[(34*4)+3] <= 1'b0;
                  spc34_inst_done         <= 0;
                  spc34_phy_pc_w          <= 0;
                end else begin
                  active_thread[(34*4)]   <= 1'b1;
                  active_thread[(34*4)+1] <= 1'b1;
                  active_thread[(34*4)+2] <= 1'b1;
                  active_thread[(34*4)+3] <= 1'b1;
                  spc34_inst_done         <= `ARIANE_CORE34.piton_pc_vld;
                  spc34_phy_pc_w          <= `ARIANE_CORE34.piton_pc;
                end
            end
    

            assign spc35_thread_id = 2'b00;
            assign spc35_rtl_pc = spc35_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(35*4)]   <= 1'b0;
                  active_thread[(35*4)+1] <= 1'b0;
                  active_thread[(35*4)+2] <= 1'b0;
                  active_thread[(35*4)+3] <= 1'b0;
                  spc35_inst_done         <= 0;
                  spc35_phy_pc_w          <= 0;
                end else begin
                  active_thread[(35*4)]   <= 1'b1;
                  active_thread[(35*4)+1] <= 1'b1;
                  active_thread[(35*4)+2] <= 1'b1;
                  active_thread[(35*4)+3] <= 1'b1;
                  spc35_inst_done         <= `ARIANE_CORE35.piton_pc_vld;
                  spc35_phy_pc_w          <= `ARIANE_CORE35.piton_pc;
                end
            end
    

            assign spc36_thread_id = 2'b00;
            assign spc36_rtl_pc = spc36_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(36*4)]   <= 1'b0;
                  active_thread[(36*4)+1] <= 1'b0;
                  active_thread[(36*4)+2] <= 1'b0;
                  active_thread[(36*4)+3] <= 1'b0;
                  spc36_inst_done         <= 0;
                  spc36_phy_pc_w          <= 0;
                end else begin
                  active_thread[(36*4)]   <= 1'b1;
                  active_thread[(36*4)+1] <= 1'b1;
                  active_thread[(36*4)+2] <= 1'b1;
                  active_thread[(36*4)+3] <= 1'b1;
                  spc36_inst_done         <= `ARIANE_CORE36.piton_pc_vld;
                  spc36_phy_pc_w          <= `ARIANE_CORE36.piton_pc;
                end
            end
    

            assign spc37_thread_id = 2'b00;
            assign spc37_rtl_pc = spc37_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(37*4)]   <= 1'b0;
                  active_thread[(37*4)+1] <= 1'b0;
                  active_thread[(37*4)+2] <= 1'b0;
                  active_thread[(37*4)+3] <= 1'b0;
                  spc37_inst_done         <= 0;
                  spc37_phy_pc_w          <= 0;
                end else begin
                  active_thread[(37*4)]   <= 1'b1;
                  active_thread[(37*4)+1] <= 1'b1;
                  active_thread[(37*4)+2] <= 1'b1;
                  active_thread[(37*4)+3] <= 1'b1;
                  spc37_inst_done         <= `ARIANE_CORE37.piton_pc_vld;
                  spc37_phy_pc_w          <= `ARIANE_CORE37.piton_pc;
                end
            end
    

            assign spc38_thread_id = 2'b00;
            assign spc38_rtl_pc = spc38_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(38*4)]   <= 1'b0;
                  active_thread[(38*4)+1] <= 1'b0;
                  active_thread[(38*4)+2] <= 1'b0;
                  active_thread[(38*4)+3] <= 1'b0;
                  spc38_inst_done         <= 0;
                  spc38_phy_pc_w          <= 0;
                end else begin
                  active_thread[(38*4)]   <= 1'b1;
                  active_thread[(38*4)+1] <= 1'b1;
                  active_thread[(38*4)+2] <= 1'b1;
                  active_thread[(38*4)+3] <= 1'b1;
                  spc38_inst_done         <= `ARIANE_CORE38.piton_pc_vld;
                  spc38_phy_pc_w          <= `ARIANE_CORE38.piton_pc;
                end
            end
    

            assign spc39_thread_id = 2'b00;
            assign spc39_rtl_pc = spc39_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(39*4)]   <= 1'b0;
                  active_thread[(39*4)+1] <= 1'b0;
                  active_thread[(39*4)+2] <= 1'b0;
                  active_thread[(39*4)+3] <= 1'b0;
                  spc39_inst_done         <= 0;
                  spc39_phy_pc_w          <= 0;
                end else begin
                  active_thread[(39*4)]   <= 1'b1;
                  active_thread[(39*4)+1] <= 1'b1;
                  active_thread[(39*4)+2] <= 1'b1;
                  active_thread[(39*4)+3] <= 1'b1;
                  spc39_inst_done         <= `ARIANE_CORE39.piton_pc_vld;
                  spc39_phy_pc_w          <= `ARIANE_CORE39.piton_pc;
                end
            end
    

            assign spc40_thread_id = 2'b00;
            assign spc40_rtl_pc = spc40_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(40*4)]   <= 1'b0;
                  active_thread[(40*4)+1] <= 1'b0;
                  active_thread[(40*4)+2] <= 1'b0;
                  active_thread[(40*4)+3] <= 1'b0;
                  spc40_inst_done         <= 0;
                  spc40_phy_pc_w          <= 0;
                end else begin
                  active_thread[(40*4)]   <= 1'b1;
                  active_thread[(40*4)+1] <= 1'b1;
                  active_thread[(40*4)+2] <= 1'b1;
                  active_thread[(40*4)+3] <= 1'b1;
                  spc40_inst_done         <= `ARIANE_CORE40.piton_pc_vld;
                  spc40_phy_pc_w          <= `ARIANE_CORE40.piton_pc;
                end
            end
    

            assign spc41_thread_id = 2'b00;
            assign spc41_rtl_pc = spc41_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(41*4)]   <= 1'b0;
                  active_thread[(41*4)+1] <= 1'b0;
                  active_thread[(41*4)+2] <= 1'b0;
                  active_thread[(41*4)+3] <= 1'b0;
                  spc41_inst_done         <= 0;
                  spc41_phy_pc_w          <= 0;
                end else begin
                  active_thread[(41*4)]   <= 1'b1;
                  active_thread[(41*4)+1] <= 1'b1;
                  active_thread[(41*4)+2] <= 1'b1;
                  active_thread[(41*4)+3] <= 1'b1;
                  spc41_inst_done         <= `ARIANE_CORE41.piton_pc_vld;
                  spc41_phy_pc_w          <= `ARIANE_CORE41.piton_pc;
                end
            end
    

            assign spc42_thread_id = 2'b00;
            assign spc42_rtl_pc = spc42_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(42*4)]   <= 1'b0;
                  active_thread[(42*4)+1] <= 1'b0;
                  active_thread[(42*4)+2] <= 1'b0;
                  active_thread[(42*4)+3] <= 1'b0;
                  spc42_inst_done         <= 0;
                  spc42_phy_pc_w          <= 0;
                end else begin
                  active_thread[(42*4)]   <= 1'b1;
                  active_thread[(42*4)+1] <= 1'b1;
                  active_thread[(42*4)+2] <= 1'b1;
                  active_thread[(42*4)+3] <= 1'b1;
                  spc42_inst_done         <= `ARIANE_CORE42.piton_pc_vld;
                  spc42_phy_pc_w          <= `ARIANE_CORE42.piton_pc;
                end
            end
    

            assign spc43_thread_id = 2'b00;
            assign spc43_rtl_pc = spc43_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(43*4)]   <= 1'b0;
                  active_thread[(43*4)+1] <= 1'b0;
                  active_thread[(43*4)+2] <= 1'b0;
                  active_thread[(43*4)+3] <= 1'b0;
                  spc43_inst_done         <= 0;
                  spc43_phy_pc_w          <= 0;
                end else begin
                  active_thread[(43*4)]   <= 1'b1;
                  active_thread[(43*4)+1] <= 1'b1;
                  active_thread[(43*4)+2] <= 1'b1;
                  active_thread[(43*4)+3] <= 1'b1;
                  spc43_inst_done         <= `ARIANE_CORE43.piton_pc_vld;
                  spc43_phy_pc_w          <= `ARIANE_CORE43.piton_pc;
                end
            end
    

            assign spc44_thread_id = 2'b00;
            assign spc44_rtl_pc = spc44_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(44*4)]   <= 1'b0;
                  active_thread[(44*4)+1] <= 1'b0;
                  active_thread[(44*4)+2] <= 1'b0;
                  active_thread[(44*4)+3] <= 1'b0;
                  spc44_inst_done         <= 0;
                  spc44_phy_pc_w          <= 0;
                end else begin
                  active_thread[(44*4)]   <= 1'b1;
                  active_thread[(44*4)+1] <= 1'b1;
                  active_thread[(44*4)+2] <= 1'b1;
                  active_thread[(44*4)+3] <= 1'b1;
                  spc44_inst_done         <= `ARIANE_CORE44.piton_pc_vld;
                  spc44_phy_pc_w          <= `ARIANE_CORE44.piton_pc;
                end
            end
    

            assign spc45_thread_id = 2'b00;
            assign spc45_rtl_pc = spc45_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(45*4)]   <= 1'b0;
                  active_thread[(45*4)+1] <= 1'b0;
                  active_thread[(45*4)+2] <= 1'b0;
                  active_thread[(45*4)+3] <= 1'b0;
                  spc45_inst_done         <= 0;
                  spc45_phy_pc_w          <= 0;
                end else begin
                  active_thread[(45*4)]   <= 1'b1;
                  active_thread[(45*4)+1] <= 1'b1;
                  active_thread[(45*4)+2] <= 1'b1;
                  active_thread[(45*4)+3] <= 1'b1;
                  spc45_inst_done         <= `ARIANE_CORE45.piton_pc_vld;
                  spc45_phy_pc_w          <= `ARIANE_CORE45.piton_pc;
                end
            end
    

            assign spc46_thread_id = 2'b00;
            assign spc46_rtl_pc = spc46_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(46*4)]   <= 1'b0;
                  active_thread[(46*4)+1] <= 1'b0;
                  active_thread[(46*4)+2] <= 1'b0;
                  active_thread[(46*4)+3] <= 1'b0;
                  spc46_inst_done         <= 0;
                  spc46_phy_pc_w          <= 0;
                end else begin
                  active_thread[(46*4)]   <= 1'b1;
                  active_thread[(46*4)+1] <= 1'b1;
                  active_thread[(46*4)+2] <= 1'b1;
                  active_thread[(46*4)+3] <= 1'b1;
                  spc46_inst_done         <= `ARIANE_CORE46.piton_pc_vld;
                  spc46_phy_pc_w          <= `ARIANE_CORE46.piton_pc;
                end
            end
    

            assign spc47_thread_id = 2'b00;
            assign spc47_rtl_pc = spc47_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(47*4)]   <= 1'b0;
                  active_thread[(47*4)+1] <= 1'b0;
                  active_thread[(47*4)+2] <= 1'b0;
                  active_thread[(47*4)+3] <= 1'b0;
                  spc47_inst_done         <= 0;
                  spc47_phy_pc_w          <= 0;
                end else begin
                  active_thread[(47*4)]   <= 1'b1;
                  active_thread[(47*4)+1] <= 1'b1;
                  active_thread[(47*4)+2] <= 1'b1;
                  active_thread[(47*4)+3] <= 1'b1;
                  spc47_inst_done         <= `ARIANE_CORE47.piton_pc_vld;
                  spc47_phy_pc_w          <= `ARIANE_CORE47.piton_pc;
                end
            end
    

            assign spc48_thread_id = 2'b00;
            assign spc48_rtl_pc = spc48_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(48*4)]   <= 1'b0;
                  active_thread[(48*4)+1] <= 1'b0;
                  active_thread[(48*4)+2] <= 1'b0;
                  active_thread[(48*4)+3] <= 1'b0;
                  spc48_inst_done         <= 0;
                  spc48_phy_pc_w          <= 0;
                end else begin
                  active_thread[(48*4)]   <= 1'b1;
                  active_thread[(48*4)+1] <= 1'b1;
                  active_thread[(48*4)+2] <= 1'b1;
                  active_thread[(48*4)+3] <= 1'b1;
                  spc48_inst_done         <= `ARIANE_CORE48.piton_pc_vld;
                  spc48_phy_pc_w          <= `ARIANE_CORE48.piton_pc;
                end
            end
    

            assign spc49_thread_id = 2'b00;
            assign spc49_rtl_pc = spc49_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(49*4)]   <= 1'b0;
                  active_thread[(49*4)+1] <= 1'b0;
                  active_thread[(49*4)+2] <= 1'b0;
                  active_thread[(49*4)+3] <= 1'b0;
                  spc49_inst_done         <= 0;
                  spc49_phy_pc_w          <= 0;
                end else begin
                  active_thread[(49*4)]   <= 1'b1;
                  active_thread[(49*4)+1] <= 1'b1;
                  active_thread[(49*4)+2] <= 1'b1;
                  active_thread[(49*4)+3] <= 1'b1;
                  spc49_inst_done         <= `ARIANE_CORE49.piton_pc_vld;
                  spc49_phy_pc_w          <= `ARIANE_CORE49.piton_pc;
                end
            end
    

            assign spc50_thread_id = 2'b00;
            assign spc50_rtl_pc = spc50_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(50*4)]   <= 1'b0;
                  active_thread[(50*4)+1] <= 1'b0;
                  active_thread[(50*4)+2] <= 1'b0;
                  active_thread[(50*4)+3] <= 1'b0;
                  spc50_inst_done         <= 0;
                  spc50_phy_pc_w          <= 0;
                end else begin
                  active_thread[(50*4)]   <= 1'b1;
                  active_thread[(50*4)+1] <= 1'b1;
                  active_thread[(50*4)+2] <= 1'b1;
                  active_thread[(50*4)+3] <= 1'b1;
                  spc50_inst_done         <= `ARIANE_CORE50.piton_pc_vld;
                  spc50_phy_pc_w          <= `ARIANE_CORE50.piton_pc;
                end
            end
    

            assign spc51_thread_id = 2'b00;
            assign spc51_rtl_pc = spc51_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(51*4)]   <= 1'b0;
                  active_thread[(51*4)+1] <= 1'b0;
                  active_thread[(51*4)+2] <= 1'b0;
                  active_thread[(51*4)+3] <= 1'b0;
                  spc51_inst_done         <= 0;
                  spc51_phy_pc_w          <= 0;
                end else begin
                  active_thread[(51*4)]   <= 1'b1;
                  active_thread[(51*4)+1] <= 1'b1;
                  active_thread[(51*4)+2] <= 1'b1;
                  active_thread[(51*4)+3] <= 1'b1;
                  spc51_inst_done         <= `ARIANE_CORE51.piton_pc_vld;
                  spc51_phy_pc_w          <= `ARIANE_CORE51.piton_pc;
                end
            end
    

            assign spc52_thread_id = 2'b00;
            assign spc52_rtl_pc = spc52_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(52*4)]   <= 1'b0;
                  active_thread[(52*4)+1] <= 1'b0;
                  active_thread[(52*4)+2] <= 1'b0;
                  active_thread[(52*4)+3] <= 1'b0;
                  spc52_inst_done         <= 0;
                  spc52_phy_pc_w          <= 0;
                end else begin
                  active_thread[(52*4)]   <= 1'b1;
                  active_thread[(52*4)+1] <= 1'b1;
                  active_thread[(52*4)+2] <= 1'b1;
                  active_thread[(52*4)+3] <= 1'b1;
                  spc52_inst_done         <= `ARIANE_CORE52.piton_pc_vld;
                  spc52_phy_pc_w          <= `ARIANE_CORE52.piton_pc;
                end
            end
    

            assign spc53_thread_id = 2'b00;
            assign spc53_rtl_pc = spc53_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(53*4)]   <= 1'b0;
                  active_thread[(53*4)+1] <= 1'b0;
                  active_thread[(53*4)+2] <= 1'b0;
                  active_thread[(53*4)+3] <= 1'b0;
                  spc53_inst_done         <= 0;
                  spc53_phy_pc_w          <= 0;
                end else begin
                  active_thread[(53*4)]   <= 1'b1;
                  active_thread[(53*4)+1] <= 1'b1;
                  active_thread[(53*4)+2] <= 1'b1;
                  active_thread[(53*4)+3] <= 1'b1;
                  spc53_inst_done         <= `ARIANE_CORE53.piton_pc_vld;
                  spc53_phy_pc_w          <= `ARIANE_CORE53.piton_pc;
                end
            end
    

            assign spc54_thread_id = 2'b00;
            assign spc54_rtl_pc = spc54_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(54*4)]   <= 1'b0;
                  active_thread[(54*4)+1] <= 1'b0;
                  active_thread[(54*4)+2] <= 1'b0;
                  active_thread[(54*4)+3] <= 1'b0;
                  spc54_inst_done         <= 0;
                  spc54_phy_pc_w          <= 0;
                end else begin
                  active_thread[(54*4)]   <= 1'b1;
                  active_thread[(54*4)+1] <= 1'b1;
                  active_thread[(54*4)+2] <= 1'b1;
                  active_thread[(54*4)+3] <= 1'b1;
                  spc54_inst_done         <= `ARIANE_CORE54.piton_pc_vld;
                  spc54_phy_pc_w          <= `ARIANE_CORE54.piton_pc;
                end
            end
    

            assign spc55_thread_id = 2'b00;
            assign spc55_rtl_pc = spc55_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(55*4)]   <= 1'b0;
                  active_thread[(55*4)+1] <= 1'b0;
                  active_thread[(55*4)+2] <= 1'b0;
                  active_thread[(55*4)+3] <= 1'b0;
                  spc55_inst_done         <= 0;
                  spc55_phy_pc_w          <= 0;
                end else begin
                  active_thread[(55*4)]   <= 1'b1;
                  active_thread[(55*4)+1] <= 1'b1;
                  active_thread[(55*4)+2] <= 1'b1;
                  active_thread[(55*4)+3] <= 1'b1;
                  spc55_inst_done         <= `ARIANE_CORE55.piton_pc_vld;
                  spc55_phy_pc_w          <= `ARIANE_CORE55.piton_pc;
                end
            end
    

            assign spc56_thread_id = 2'b00;
            assign spc56_rtl_pc = spc56_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(56*4)]   <= 1'b0;
                  active_thread[(56*4)+1] <= 1'b0;
                  active_thread[(56*4)+2] <= 1'b0;
                  active_thread[(56*4)+3] <= 1'b0;
                  spc56_inst_done         <= 0;
                  spc56_phy_pc_w          <= 0;
                end else begin
                  active_thread[(56*4)]   <= 1'b1;
                  active_thread[(56*4)+1] <= 1'b1;
                  active_thread[(56*4)+2] <= 1'b1;
                  active_thread[(56*4)+3] <= 1'b1;
                  spc56_inst_done         <= `ARIANE_CORE56.piton_pc_vld;
                  spc56_phy_pc_w          <= `ARIANE_CORE56.piton_pc;
                end
            end
    

            assign spc57_thread_id = 2'b00;
            assign spc57_rtl_pc = spc57_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(57*4)]   <= 1'b0;
                  active_thread[(57*4)+1] <= 1'b0;
                  active_thread[(57*4)+2] <= 1'b0;
                  active_thread[(57*4)+3] <= 1'b0;
                  spc57_inst_done         <= 0;
                  spc57_phy_pc_w          <= 0;
                end else begin
                  active_thread[(57*4)]   <= 1'b1;
                  active_thread[(57*4)+1] <= 1'b1;
                  active_thread[(57*4)+2] <= 1'b1;
                  active_thread[(57*4)+3] <= 1'b1;
                  spc57_inst_done         <= `ARIANE_CORE57.piton_pc_vld;
                  spc57_phy_pc_w          <= `ARIANE_CORE57.piton_pc;
                end
            end
    

            assign spc58_thread_id = 2'b00;
            assign spc58_rtl_pc = spc58_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(58*4)]   <= 1'b0;
                  active_thread[(58*4)+1] <= 1'b0;
                  active_thread[(58*4)+2] <= 1'b0;
                  active_thread[(58*4)+3] <= 1'b0;
                  spc58_inst_done         <= 0;
                  spc58_phy_pc_w          <= 0;
                end else begin
                  active_thread[(58*4)]   <= 1'b1;
                  active_thread[(58*4)+1] <= 1'b1;
                  active_thread[(58*4)+2] <= 1'b1;
                  active_thread[(58*4)+3] <= 1'b1;
                  spc58_inst_done         <= `ARIANE_CORE58.piton_pc_vld;
                  spc58_phy_pc_w          <= `ARIANE_CORE58.piton_pc;
                end
            end
    

            assign spc59_thread_id = 2'b00;
            assign spc59_rtl_pc = spc59_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(59*4)]   <= 1'b0;
                  active_thread[(59*4)+1] <= 1'b0;
                  active_thread[(59*4)+2] <= 1'b0;
                  active_thread[(59*4)+3] <= 1'b0;
                  spc59_inst_done         <= 0;
                  spc59_phy_pc_w          <= 0;
                end else begin
                  active_thread[(59*4)]   <= 1'b1;
                  active_thread[(59*4)+1] <= 1'b1;
                  active_thread[(59*4)+2] <= 1'b1;
                  active_thread[(59*4)+3] <= 1'b1;
                  spc59_inst_done         <= `ARIANE_CORE59.piton_pc_vld;
                  spc59_phy_pc_w          <= `ARIANE_CORE59.piton_pc;
                end
            end
    

            assign spc60_thread_id = 2'b00;
            assign spc60_rtl_pc = spc60_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(60*4)]   <= 1'b0;
                  active_thread[(60*4)+1] <= 1'b0;
                  active_thread[(60*4)+2] <= 1'b0;
                  active_thread[(60*4)+3] <= 1'b0;
                  spc60_inst_done         <= 0;
                  spc60_phy_pc_w          <= 0;
                end else begin
                  active_thread[(60*4)]   <= 1'b1;
                  active_thread[(60*4)+1] <= 1'b1;
                  active_thread[(60*4)+2] <= 1'b1;
                  active_thread[(60*4)+3] <= 1'b1;
                  spc60_inst_done         <= `ARIANE_CORE60.piton_pc_vld;
                  spc60_phy_pc_w          <= `ARIANE_CORE60.piton_pc;
                end
            end
    

            assign spc61_thread_id = 2'b00;
            assign spc61_rtl_pc = spc61_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(61*4)]   <= 1'b0;
                  active_thread[(61*4)+1] <= 1'b0;
                  active_thread[(61*4)+2] <= 1'b0;
                  active_thread[(61*4)+3] <= 1'b0;
                  spc61_inst_done         <= 0;
                  spc61_phy_pc_w          <= 0;
                end else begin
                  active_thread[(61*4)]   <= 1'b1;
                  active_thread[(61*4)+1] <= 1'b1;
                  active_thread[(61*4)+2] <= 1'b1;
                  active_thread[(61*4)+3] <= 1'b1;
                  spc61_inst_done         <= `ARIANE_CORE61.piton_pc_vld;
                  spc61_phy_pc_w          <= `ARIANE_CORE61.piton_pc;
                end
            end
    

            assign spc62_thread_id = 2'b00;
            assign spc62_rtl_pc = spc62_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(62*4)]   <= 1'b0;
                  active_thread[(62*4)+1] <= 1'b0;
                  active_thread[(62*4)+2] <= 1'b0;
                  active_thread[(62*4)+3] <= 1'b0;
                  spc62_inst_done         <= 0;
                  spc62_phy_pc_w          <= 0;
                end else begin
                  active_thread[(62*4)]   <= 1'b1;
                  active_thread[(62*4)+1] <= 1'b1;
                  active_thread[(62*4)+2] <= 1'b1;
                  active_thread[(62*4)+3] <= 1'b1;
                  spc62_inst_done         <= `ARIANE_CORE62.piton_pc_vld;
                  spc62_phy_pc_w          <= `ARIANE_CORE62.piton_pc;
                end
            end
    

            assign spc63_thread_id = 2'b00;
            assign spc63_rtl_pc = spc63_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(63*4)]   <= 1'b0;
                  active_thread[(63*4)+1] <= 1'b0;
                  active_thread[(63*4)+2] <= 1'b0;
                  active_thread[(63*4)+3] <= 1'b0;
                  spc63_inst_done         <= 0;
                  spc63_phy_pc_w          <= 0;
                end else begin
                  active_thread[(63*4)]   <= 1'b1;
                  active_thread[(63*4)+1] <= 1'b1;
                  active_thread[(63*4)+2] <= 1'b1;
                  active_thread[(63*4)+3] <= 1'b1;
                  spc63_inst_done         <= `ARIANE_CORE63.piton_pc_vld;
                  spc63_phy_pc_w          <= `ARIANE_CORE63.piton_pc;
                end
            end
    

            assign spc64_thread_id = 2'b00;
            assign spc64_rtl_pc = spc64_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(64*4)]   <= 1'b0;
                  active_thread[(64*4)+1] <= 1'b0;
                  active_thread[(64*4)+2] <= 1'b0;
                  active_thread[(64*4)+3] <= 1'b0;
                  spc64_inst_done         <= 0;
                  spc64_phy_pc_w          <= 0;
                end else begin
                  active_thread[(64*4)]   <= 1'b1;
                  active_thread[(64*4)+1] <= 1'b1;
                  active_thread[(64*4)+2] <= 1'b1;
                  active_thread[(64*4)+3] <= 1'b1;
                  spc64_inst_done         <= `ARIANE_CORE64.piton_pc_vld;
                  spc64_phy_pc_w          <= `ARIANE_CORE64.piton_pc;
                end
            end
    

            assign spc65_thread_id = 2'b00;
            assign spc65_rtl_pc = spc65_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(65*4)]   <= 1'b0;
                  active_thread[(65*4)+1] <= 1'b0;
                  active_thread[(65*4)+2] <= 1'b0;
                  active_thread[(65*4)+3] <= 1'b0;
                  spc65_inst_done         <= 0;
                  spc65_phy_pc_w          <= 0;
                end else begin
                  active_thread[(65*4)]   <= 1'b1;
                  active_thread[(65*4)+1] <= 1'b1;
                  active_thread[(65*4)+2] <= 1'b1;
                  active_thread[(65*4)+3] <= 1'b1;
                  spc65_inst_done         <= `ARIANE_CORE65.piton_pc_vld;
                  spc65_phy_pc_w          <= `ARIANE_CORE65.piton_pc;
                end
            end
    

            assign spc66_thread_id = 2'b00;
            assign spc66_rtl_pc = spc66_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(66*4)]   <= 1'b0;
                  active_thread[(66*4)+1] <= 1'b0;
                  active_thread[(66*4)+2] <= 1'b0;
                  active_thread[(66*4)+3] <= 1'b0;
                  spc66_inst_done         <= 0;
                  spc66_phy_pc_w          <= 0;
                end else begin
                  active_thread[(66*4)]   <= 1'b1;
                  active_thread[(66*4)+1] <= 1'b1;
                  active_thread[(66*4)+2] <= 1'b1;
                  active_thread[(66*4)+3] <= 1'b1;
                  spc66_inst_done         <= `ARIANE_CORE66.piton_pc_vld;
                  spc66_phy_pc_w          <= `ARIANE_CORE66.piton_pc;
                end
            end
    

            assign spc67_thread_id = 2'b00;
            assign spc67_rtl_pc = spc67_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(67*4)]   <= 1'b0;
                  active_thread[(67*4)+1] <= 1'b0;
                  active_thread[(67*4)+2] <= 1'b0;
                  active_thread[(67*4)+3] <= 1'b0;
                  spc67_inst_done         <= 0;
                  spc67_phy_pc_w          <= 0;
                end else begin
                  active_thread[(67*4)]   <= 1'b1;
                  active_thread[(67*4)+1] <= 1'b1;
                  active_thread[(67*4)+2] <= 1'b1;
                  active_thread[(67*4)+3] <= 1'b1;
                  spc67_inst_done         <= `ARIANE_CORE67.piton_pc_vld;
                  spc67_phy_pc_w          <= `ARIANE_CORE67.piton_pc;
                end
            end
    

            assign spc68_thread_id = 2'b00;
            assign spc68_rtl_pc = spc68_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(68*4)]   <= 1'b0;
                  active_thread[(68*4)+1] <= 1'b0;
                  active_thread[(68*4)+2] <= 1'b0;
                  active_thread[(68*4)+3] <= 1'b0;
                  spc68_inst_done         <= 0;
                  spc68_phy_pc_w          <= 0;
                end else begin
                  active_thread[(68*4)]   <= 1'b1;
                  active_thread[(68*4)+1] <= 1'b1;
                  active_thread[(68*4)+2] <= 1'b1;
                  active_thread[(68*4)+3] <= 1'b1;
                  spc68_inst_done         <= `ARIANE_CORE68.piton_pc_vld;
                  spc68_phy_pc_w          <= `ARIANE_CORE68.piton_pc;
                end
            end
    

            assign spc69_thread_id = 2'b00;
            assign spc69_rtl_pc = spc69_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(69*4)]   <= 1'b0;
                  active_thread[(69*4)+1] <= 1'b0;
                  active_thread[(69*4)+2] <= 1'b0;
                  active_thread[(69*4)+3] <= 1'b0;
                  spc69_inst_done         <= 0;
                  spc69_phy_pc_w          <= 0;
                end else begin
                  active_thread[(69*4)]   <= 1'b1;
                  active_thread[(69*4)+1] <= 1'b1;
                  active_thread[(69*4)+2] <= 1'b1;
                  active_thread[(69*4)+3] <= 1'b1;
                  spc69_inst_done         <= `ARIANE_CORE69.piton_pc_vld;
                  spc69_phy_pc_w          <= `ARIANE_CORE69.piton_pc;
                end
            end
    

            assign spc70_thread_id = 2'b00;
            assign spc70_rtl_pc = spc70_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(70*4)]   <= 1'b0;
                  active_thread[(70*4)+1] <= 1'b0;
                  active_thread[(70*4)+2] <= 1'b0;
                  active_thread[(70*4)+3] <= 1'b0;
                  spc70_inst_done         <= 0;
                  spc70_phy_pc_w          <= 0;
                end else begin
                  active_thread[(70*4)]   <= 1'b1;
                  active_thread[(70*4)+1] <= 1'b1;
                  active_thread[(70*4)+2] <= 1'b1;
                  active_thread[(70*4)+3] <= 1'b1;
                  spc70_inst_done         <= `ARIANE_CORE70.piton_pc_vld;
                  spc70_phy_pc_w          <= `ARIANE_CORE70.piton_pc;
                end
            end
    

            assign spc71_thread_id = 2'b00;
            assign spc71_rtl_pc = spc71_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(71*4)]   <= 1'b0;
                  active_thread[(71*4)+1] <= 1'b0;
                  active_thread[(71*4)+2] <= 1'b0;
                  active_thread[(71*4)+3] <= 1'b0;
                  spc71_inst_done         <= 0;
                  spc71_phy_pc_w          <= 0;
                end else begin
                  active_thread[(71*4)]   <= 1'b1;
                  active_thread[(71*4)+1] <= 1'b1;
                  active_thread[(71*4)+2] <= 1'b1;
                  active_thread[(71*4)+3] <= 1'b1;
                  spc71_inst_done         <= `ARIANE_CORE71.piton_pc_vld;
                  spc71_phy_pc_w          <= `ARIANE_CORE71.piton_pc;
                end
            end
    

            assign spc72_thread_id = 2'b00;
            assign spc72_rtl_pc = spc72_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(72*4)]   <= 1'b0;
                  active_thread[(72*4)+1] <= 1'b0;
                  active_thread[(72*4)+2] <= 1'b0;
                  active_thread[(72*4)+3] <= 1'b0;
                  spc72_inst_done         <= 0;
                  spc72_phy_pc_w          <= 0;
                end else begin
                  active_thread[(72*4)]   <= 1'b1;
                  active_thread[(72*4)+1] <= 1'b1;
                  active_thread[(72*4)+2] <= 1'b1;
                  active_thread[(72*4)+3] <= 1'b1;
                  spc72_inst_done         <= `ARIANE_CORE72.piton_pc_vld;
                  spc72_phy_pc_w          <= `ARIANE_CORE72.piton_pc;
                end
            end
    

            assign spc73_thread_id = 2'b00;
            assign spc73_rtl_pc = spc73_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(73*4)]   <= 1'b0;
                  active_thread[(73*4)+1] <= 1'b0;
                  active_thread[(73*4)+2] <= 1'b0;
                  active_thread[(73*4)+3] <= 1'b0;
                  spc73_inst_done         <= 0;
                  spc73_phy_pc_w          <= 0;
                end else begin
                  active_thread[(73*4)]   <= 1'b1;
                  active_thread[(73*4)+1] <= 1'b1;
                  active_thread[(73*4)+2] <= 1'b1;
                  active_thread[(73*4)+3] <= 1'b1;
                  spc73_inst_done         <= `ARIANE_CORE73.piton_pc_vld;
                  spc73_phy_pc_w          <= `ARIANE_CORE73.piton_pc;
                end
            end
    

            assign spc74_thread_id = 2'b00;
            assign spc74_rtl_pc = spc74_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(74*4)]   <= 1'b0;
                  active_thread[(74*4)+1] <= 1'b0;
                  active_thread[(74*4)+2] <= 1'b0;
                  active_thread[(74*4)+3] <= 1'b0;
                  spc74_inst_done         <= 0;
                  spc74_phy_pc_w          <= 0;
                end else begin
                  active_thread[(74*4)]   <= 1'b1;
                  active_thread[(74*4)+1] <= 1'b1;
                  active_thread[(74*4)+2] <= 1'b1;
                  active_thread[(74*4)+3] <= 1'b1;
                  spc74_inst_done         <= `ARIANE_CORE74.piton_pc_vld;
                  spc74_phy_pc_w          <= `ARIANE_CORE74.piton_pc;
                end
            end
    

            assign spc75_thread_id = 2'b00;
            assign spc75_rtl_pc = spc75_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(75*4)]   <= 1'b0;
                  active_thread[(75*4)+1] <= 1'b0;
                  active_thread[(75*4)+2] <= 1'b0;
                  active_thread[(75*4)+3] <= 1'b0;
                  spc75_inst_done         <= 0;
                  spc75_phy_pc_w          <= 0;
                end else begin
                  active_thread[(75*4)]   <= 1'b1;
                  active_thread[(75*4)+1] <= 1'b1;
                  active_thread[(75*4)+2] <= 1'b1;
                  active_thread[(75*4)+3] <= 1'b1;
                  spc75_inst_done         <= `ARIANE_CORE75.piton_pc_vld;
                  spc75_phy_pc_w          <= `ARIANE_CORE75.piton_pc;
                end
            end
    

            assign spc76_thread_id = 2'b00;
            assign spc76_rtl_pc = spc76_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(76*4)]   <= 1'b0;
                  active_thread[(76*4)+1] <= 1'b0;
                  active_thread[(76*4)+2] <= 1'b0;
                  active_thread[(76*4)+3] <= 1'b0;
                  spc76_inst_done         <= 0;
                  spc76_phy_pc_w          <= 0;
                end else begin
                  active_thread[(76*4)]   <= 1'b1;
                  active_thread[(76*4)+1] <= 1'b1;
                  active_thread[(76*4)+2] <= 1'b1;
                  active_thread[(76*4)+3] <= 1'b1;
                  spc76_inst_done         <= `ARIANE_CORE76.piton_pc_vld;
                  spc76_phy_pc_w          <= `ARIANE_CORE76.piton_pc;
                end
            end
    

            assign spc77_thread_id = 2'b00;
            assign spc77_rtl_pc = spc77_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(77*4)]   <= 1'b0;
                  active_thread[(77*4)+1] <= 1'b0;
                  active_thread[(77*4)+2] <= 1'b0;
                  active_thread[(77*4)+3] <= 1'b0;
                  spc77_inst_done         <= 0;
                  spc77_phy_pc_w          <= 0;
                end else begin
                  active_thread[(77*4)]   <= 1'b1;
                  active_thread[(77*4)+1] <= 1'b1;
                  active_thread[(77*4)+2] <= 1'b1;
                  active_thread[(77*4)+3] <= 1'b1;
                  spc77_inst_done         <= `ARIANE_CORE77.piton_pc_vld;
                  spc77_phy_pc_w          <= `ARIANE_CORE77.piton_pc;
                end
            end
    

            assign spc78_thread_id = 2'b00;
            assign spc78_rtl_pc = spc78_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(78*4)]   <= 1'b0;
                  active_thread[(78*4)+1] <= 1'b0;
                  active_thread[(78*4)+2] <= 1'b0;
                  active_thread[(78*4)+3] <= 1'b0;
                  spc78_inst_done         <= 0;
                  spc78_phy_pc_w          <= 0;
                end else begin
                  active_thread[(78*4)]   <= 1'b1;
                  active_thread[(78*4)+1] <= 1'b1;
                  active_thread[(78*4)+2] <= 1'b1;
                  active_thread[(78*4)+3] <= 1'b1;
                  spc78_inst_done         <= `ARIANE_CORE78.piton_pc_vld;
                  spc78_phy_pc_w          <= `ARIANE_CORE78.piton_pc;
                end
            end
    

            assign spc79_thread_id = 2'b00;
            assign spc79_rtl_pc = spc79_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(79*4)]   <= 1'b0;
                  active_thread[(79*4)+1] <= 1'b0;
                  active_thread[(79*4)+2] <= 1'b0;
                  active_thread[(79*4)+3] <= 1'b0;
                  spc79_inst_done         <= 0;
                  spc79_phy_pc_w          <= 0;
                end else begin
                  active_thread[(79*4)]   <= 1'b1;
                  active_thread[(79*4)+1] <= 1'b1;
                  active_thread[(79*4)+2] <= 1'b1;
                  active_thread[(79*4)+3] <= 1'b1;
                  spc79_inst_done         <= `ARIANE_CORE79.piton_pc_vld;
                  spc79_phy_pc_w          <= `ARIANE_CORE79.piton_pc;
                end
            end
    

            assign spc80_thread_id = 2'b00;
            assign spc80_rtl_pc = spc80_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(80*4)]   <= 1'b0;
                  active_thread[(80*4)+1] <= 1'b0;
                  active_thread[(80*4)+2] <= 1'b0;
                  active_thread[(80*4)+3] <= 1'b0;
                  spc80_inst_done         <= 0;
                  spc80_phy_pc_w          <= 0;
                end else begin
                  active_thread[(80*4)]   <= 1'b1;
                  active_thread[(80*4)+1] <= 1'b1;
                  active_thread[(80*4)+2] <= 1'b1;
                  active_thread[(80*4)+3] <= 1'b1;
                  spc80_inst_done         <= `ARIANE_CORE80.piton_pc_vld;
                  spc80_phy_pc_w          <= `ARIANE_CORE80.piton_pc;
                end
            end
    

            assign spc81_thread_id = 2'b00;
            assign spc81_rtl_pc = spc81_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(81*4)]   <= 1'b0;
                  active_thread[(81*4)+1] <= 1'b0;
                  active_thread[(81*4)+2] <= 1'b0;
                  active_thread[(81*4)+3] <= 1'b0;
                  spc81_inst_done         <= 0;
                  spc81_phy_pc_w          <= 0;
                end else begin
                  active_thread[(81*4)]   <= 1'b1;
                  active_thread[(81*4)+1] <= 1'b1;
                  active_thread[(81*4)+2] <= 1'b1;
                  active_thread[(81*4)+3] <= 1'b1;
                  spc81_inst_done         <= `ARIANE_CORE81.piton_pc_vld;
                  spc81_phy_pc_w          <= `ARIANE_CORE81.piton_pc;
                end
            end
    

            assign spc82_thread_id = 2'b00;
            assign spc82_rtl_pc = spc82_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(82*4)]   <= 1'b0;
                  active_thread[(82*4)+1] <= 1'b0;
                  active_thread[(82*4)+2] <= 1'b0;
                  active_thread[(82*4)+3] <= 1'b0;
                  spc82_inst_done         <= 0;
                  spc82_phy_pc_w          <= 0;
                end else begin
                  active_thread[(82*4)]   <= 1'b1;
                  active_thread[(82*4)+1] <= 1'b1;
                  active_thread[(82*4)+2] <= 1'b1;
                  active_thread[(82*4)+3] <= 1'b1;
                  spc82_inst_done         <= `ARIANE_CORE82.piton_pc_vld;
                  spc82_phy_pc_w          <= `ARIANE_CORE82.piton_pc;
                end
            end
    

            assign spc83_thread_id = 2'b00;
            assign spc83_rtl_pc = spc83_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(83*4)]   <= 1'b0;
                  active_thread[(83*4)+1] <= 1'b0;
                  active_thread[(83*4)+2] <= 1'b0;
                  active_thread[(83*4)+3] <= 1'b0;
                  spc83_inst_done         <= 0;
                  spc83_phy_pc_w          <= 0;
                end else begin
                  active_thread[(83*4)]   <= 1'b1;
                  active_thread[(83*4)+1] <= 1'b1;
                  active_thread[(83*4)+2] <= 1'b1;
                  active_thread[(83*4)+3] <= 1'b1;
                  spc83_inst_done         <= `ARIANE_CORE83.piton_pc_vld;
                  spc83_phy_pc_w          <= `ARIANE_CORE83.piton_pc;
                end
            end
    

            assign spc84_thread_id = 2'b00;
            assign spc84_rtl_pc = spc84_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(84*4)]   <= 1'b0;
                  active_thread[(84*4)+1] <= 1'b0;
                  active_thread[(84*4)+2] <= 1'b0;
                  active_thread[(84*4)+3] <= 1'b0;
                  spc84_inst_done         <= 0;
                  spc84_phy_pc_w          <= 0;
                end else begin
                  active_thread[(84*4)]   <= 1'b1;
                  active_thread[(84*4)+1] <= 1'b1;
                  active_thread[(84*4)+2] <= 1'b1;
                  active_thread[(84*4)+3] <= 1'b1;
                  spc84_inst_done         <= `ARIANE_CORE84.piton_pc_vld;
                  spc84_phy_pc_w          <= `ARIANE_CORE84.piton_pc;
                end
            end
    

            assign spc85_thread_id = 2'b00;
            assign spc85_rtl_pc = spc85_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(85*4)]   <= 1'b0;
                  active_thread[(85*4)+1] <= 1'b0;
                  active_thread[(85*4)+2] <= 1'b0;
                  active_thread[(85*4)+3] <= 1'b0;
                  spc85_inst_done         <= 0;
                  spc85_phy_pc_w          <= 0;
                end else begin
                  active_thread[(85*4)]   <= 1'b1;
                  active_thread[(85*4)+1] <= 1'b1;
                  active_thread[(85*4)+2] <= 1'b1;
                  active_thread[(85*4)+3] <= 1'b1;
                  spc85_inst_done         <= `ARIANE_CORE85.piton_pc_vld;
                  spc85_phy_pc_w          <= `ARIANE_CORE85.piton_pc;
                end
            end
    

            assign spc86_thread_id = 2'b00;
            assign spc86_rtl_pc = spc86_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(86*4)]   <= 1'b0;
                  active_thread[(86*4)+1] <= 1'b0;
                  active_thread[(86*4)+2] <= 1'b0;
                  active_thread[(86*4)+3] <= 1'b0;
                  spc86_inst_done         <= 0;
                  spc86_phy_pc_w          <= 0;
                end else begin
                  active_thread[(86*4)]   <= 1'b1;
                  active_thread[(86*4)+1] <= 1'b1;
                  active_thread[(86*4)+2] <= 1'b1;
                  active_thread[(86*4)+3] <= 1'b1;
                  spc86_inst_done         <= `ARIANE_CORE86.piton_pc_vld;
                  spc86_phy_pc_w          <= `ARIANE_CORE86.piton_pc;
                end
            end
    

            assign spc87_thread_id = 2'b00;
            assign spc87_rtl_pc = spc87_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(87*4)]   <= 1'b0;
                  active_thread[(87*4)+1] <= 1'b0;
                  active_thread[(87*4)+2] <= 1'b0;
                  active_thread[(87*4)+3] <= 1'b0;
                  spc87_inst_done         <= 0;
                  spc87_phy_pc_w          <= 0;
                end else begin
                  active_thread[(87*4)]   <= 1'b1;
                  active_thread[(87*4)+1] <= 1'b1;
                  active_thread[(87*4)+2] <= 1'b1;
                  active_thread[(87*4)+3] <= 1'b1;
                  spc87_inst_done         <= `ARIANE_CORE87.piton_pc_vld;
                  spc87_phy_pc_w          <= `ARIANE_CORE87.piton_pc;
                end
            end
    

            assign spc88_thread_id = 2'b00;
            assign spc88_rtl_pc = spc88_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(88*4)]   <= 1'b0;
                  active_thread[(88*4)+1] <= 1'b0;
                  active_thread[(88*4)+2] <= 1'b0;
                  active_thread[(88*4)+3] <= 1'b0;
                  spc88_inst_done         <= 0;
                  spc88_phy_pc_w          <= 0;
                end else begin
                  active_thread[(88*4)]   <= 1'b1;
                  active_thread[(88*4)+1] <= 1'b1;
                  active_thread[(88*4)+2] <= 1'b1;
                  active_thread[(88*4)+3] <= 1'b1;
                  spc88_inst_done         <= `ARIANE_CORE88.piton_pc_vld;
                  spc88_phy_pc_w          <= `ARIANE_CORE88.piton_pc;
                end
            end
    

            assign spc89_thread_id = 2'b00;
            assign spc89_rtl_pc = spc89_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(89*4)]   <= 1'b0;
                  active_thread[(89*4)+1] <= 1'b0;
                  active_thread[(89*4)+2] <= 1'b0;
                  active_thread[(89*4)+3] <= 1'b0;
                  spc89_inst_done         <= 0;
                  spc89_phy_pc_w          <= 0;
                end else begin
                  active_thread[(89*4)]   <= 1'b1;
                  active_thread[(89*4)+1] <= 1'b1;
                  active_thread[(89*4)+2] <= 1'b1;
                  active_thread[(89*4)+3] <= 1'b1;
                  spc89_inst_done         <= `ARIANE_CORE89.piton_pc_vld;
                  spc89_phy_pc_w          <= `ARIANE_CORE89.piton_pc;
                end
            end
    

            assign spc90_thread_id = 2'b00;
            assign spc90_rtl_pc = spc90_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(90*4)]   <= 1'b0;
                  active_thread[(90*4)+1] <= 1'b0;
                  active_thread[(90*4)+2] <= 1'b0;
                  active_thread[(90*4)+3] <= 1'b0;
                  spc90_inst_done         <= 0;
                  spc90_phy_pc_w          <= 0;
                end else begin
                  active_thread[(90*4)]   <= 1'b1;
                  active_thread[(90*4)+1] <= 1'b1;
                  active_thread[(90*4)+2] <= 1'b1;
                  active_thread[(90*4)+3] <= 1'b1;
                  spc90_inst_done         <= `ARIANE_CORE90.piton_pc_vld;
                  spc90_phy_pc_w          <= `ARIANE_CORE90.piton_pc;
                end
            end
    

            assign spc91_thread_id = 2'b00;
            assign spc91_rtl_pc = spc91_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(91*4)]   <= 1'b0;
                  active_thread[(91*4)+1] <= 1'b0;
                  active_thread[(91*4)+2] <= 1'b0;
                  active_thread[(91*4)+3] <= 1'b0;
                  spc91_inst_done         <= 0;
                  spc91_phy_pc_w          <= 0;
                end else begin
                  active_thread[(91*4)]   <= 1'b1;
                  active_thread[(91*4)+1] <= 1'b1;
                  active_thread[(91*4)+2] <= 1'b1;
                  active_thread[(91*4)+3] <= 1'b1;
                  spc91_inst_done         <= `ARIANE_CORE91.piton_pc_vld;
                  spc91_phy_pc_w          <= `ARIANE_CORE91.piton_pc;
                end
            end
    

            assign spc92_thread_id = 2'b00;
            assign spc92_rtl_pc = spc92_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(92*4)]   <= 1'b0;
                  active_thread[(92*4)+1] <= 1'b0;
                  active_thread[(92*4)+2] <= 1'b0;
                  active_thread[(92*4)+3] <= 1'b0;
                  spc92_inst_done         <= 0;
                  spc92_phy_pc_w          <= 0;
                end else begin
                  active_thread[(92*4)]   <= 1'b1;
                  active_thread[(92*4)+1] <= 1'b1;
                  active_thread[(92*4)+2] <= 1'b1;
                  active_thread[(92*4)+3] <= 1'b1;
                  spc92_inst_done         <= `ARIANE_CORE92.piton_pc_vld;
                  spc92_phy_pc_w          <= `ARIANE_CORE92.piton_pc;
                end
            end
    

            assign spc93_thread_id = 2'b00;
            assign spc93_rtl_pc = spc93_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(93*4)]   <= 1'b0;
                  active_thread[(93*4)+1] <= 1'b0;
                  active_thread[(93*4)+2] <= 1'b0;
                  active_thread[(93*4)+3] <= 1'b0;
                  spc93_inst_done         <= 0;
                  spc93_phy_pc_w          <= 0;
                end else begin
                  active_thread[(93*4)]   <= 1'b1;
                  active_thread[(93*4)+1] <= 1'b1;
                  active_thread[(93*4)+2] <= 1'b1;
                  active_thread[(93*4)+3] <= 1'b1;
                  spc93_inst_done         <= `ARIANE_CORE93.piton_pc_vld;
                  spc93_phy_pc_w          <= `ARIANE_CORE93.piton_pc;
                end
            end
    

            assign spc94_thread_id = 2'b00;
            assign spc94_rtl_pc = spc94_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(94*4)]   <= 1'b0;
                  active_thread[(94*4)+1] <= 1'b0;
                  active_thread[(94*4)+2] <= 1'b0;
                  active_thread[(94*4)+3] <= 1'b0;
                  spc94_inst_done         <= 0;
                  spc94_phy_pc_w          <= 0;
                end else begin
                  active_thread[(94*4)]   <= 1'b1;
                  active_thread[(94*4)+1] <= 1'b1;
                  active_thread[(94*4)+2] <= 1'b1;
                  active_thread[(94*4)+3] <= 1'b1;
                  spc94_inst_done         <= `ARIANE_CORE94.piton_pc_vld;
                  spc94_phy_pc_w          <= `ARIANE_CORE94.piton_pc;
                end
            end
    

            assign spc95_thread_id = 2'b00;
            assign spc95_rtl_pc = spc95_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(95*4)]   <= 1'b0;
                  active_thread[(95*4)+1] <= 1'b0;
                  active_thread[(95*4)+2] <= 1'b0;
                  active_thread[(95*4)+3] <= 1'b0;
                  spc95_inst_done         <= 0;
                  spc95_phy_pc_w          <= 0;
                end else begin
                  active_thread[(95*4)]   <= 1'b1;
                  active_thread[(95*4)+1] <= 1'b1;
                  active_thread[(95*4)+2] <= 1'b1;
                  active_thread[(95*4)+3] <= 1'b1;
                  spc95_inst_done         <= `ARIANE_CORE95.piton_pc_vld;
                  spc95_phy_pc_w          <= `ARIANE_CORE95.piton_pc;
                end
            end
    

            assign spc96_thread_id = 2'b00;
            assign spc96_rtl_pc = spc96_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(96*4)]   <= 1'b0;
                  active_thread[(96*4)+1] <= 1'b0;
                  active_thread[(96*4)+2] <= 1'b0;
                  active_thread[(96*4)+3] <= 1'b0;
                  spc96_inst_done         <= 0;
                  spc96_phy_pc_w          <= 0;
                end else begin
                  active_thread[(96*4)]   <= 1'b1;
                  active_thread[(96*4)+1] <= 1'b1;
                  active_thread[(96*4)+2] <= 1'b1;
                  active_thread[(96*4)+3] <= 1'b1;
                  spc96_inst_done         <= `ARIANE_CORE96.piton_pc_vld;
                  spc96_phy_pc_w          <= `ARIANE_CORE96.piton_pc;
                end
            end
    

            assign spc97_thread_id = 2'b00;
            assign spc97_rtl_pc = spc97_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(97*4)]   <= 1'b0;
                  active_thread[(97*4)+1] <= 1'b0;
                  active_thread[(97*4)+2] <= 1'b0;
                  active_thread[(97*4)+3] <= 1'b0;
                  spc97_inst_done         <= 0;
                  spc97_phy_pc_w          <= 0;
                end else begin
                  active_thread[(97*4)]   <= 1'b1;
                  active_thread[(97*4)+1] <= 1'b1;
                  active_thread[(97*4)+2] <= 1'b1;
                  active_thread[(97*4)+3] <= 1'b1;
                  spc97_inst_done         <= `ARIANE_CORE97.piton_pc_vld;
                  spc97_phy_pc_w          <= `ARIANE_CORE97.piton_pc;
                end
            end
    

            assign spc98_thread_id = 2'b00;
            assign spc98_rtl_pc = spc98_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(98*4)]   <= 1'b0;
                  active_thread[(98*4)+1] <= 1'b0;
                  active_thread[(98*4)+2] <= 1'b0;
                  active_thread[(98*4)+3] <= 1'b0;
                  spc98_inst_done         <= 0;
                  spc98_phy_pc_w          <= 0;
                end else begin
                  active_thread[(98*4)]   <= 1'b1;
                  active_thread[(98*4)+1] <= 1'b1;
                  active_thread[(98*4)+2] <= 1'b1;
                  active_thread[(98*4)+3] <= 1'b1;
                  spc98_inst_done         <= `ARIANE_CORE98.piton_pc_vld;
                  spc98_phy_pc_w          <= `ARIANE_CORE98.piton_pc;
                end
            end
    

            assign spc99_thread_id = 2'b00;
            assign spc99_rtl_pc = spc99_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(99*4)]   <= 1'b0;
                  active_thread[(99*4)+1] <= 1'b0;
                  active_thread[(99*4)+2] <= 1'b0;
                  active_thread[(99*4)+3] <= 1'b0;
                  spc99_inst_done         <= 0;
                  spc99_phy_pc_w          <= 0;
                end else begin
                  active_thread[(99*4)]   <= 1'b1;
                  active_thread[(99*4)+1] <= 1'b1;
                  active_thread[(99*4)+2] <= 1'b1;
                  active_thread[(99*4)+3] <= 1'b1;
                  spc99_inst_done         <= `ARIANE_CORE99.piton_pc_vld;
                  spc99_phy_pc_w          <= `ARIANE_CORE99.piton_pc;
                end
            end
    

            assign spc100_thread_id = 2'b00;
            assign spc100_rtl_pc = spc100_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(100*4)]   <= 1'b0;
                  active_thread[(100*4)+1] <= 1'b0;
                  active_thread[(100*4)+2] <= 1'b0;
                  active_thread[(100*4)+3] <= 1'b0;
                  spc100_inst_done         <= 0;
                  spc100_phy_pc_w          <= 0;
                end else begin
                  active_thread[(100*4)]   <= 1'b1;
                  active_thread[(100*4)+1] <= 1'b1;
                  active_thread[(100*4)+2] <= 1'b1;
                  active_thread[(100*4)+3] <= 1'b1;
                  spc100_inst_done         <= `ARIANE_CORE100.piton_pc_vld;
                  spc100_phy_pc_w          <= `ARIANE_CORE100.piton_pc;
                end
            end
    

            assign spc101_thread_id = 2'b00;
            assign spc101_rtl_pc = spc101_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(101*4)]   <= 1'b0;
                  active_thread[(101*4)+1] <= 1'b0;
                  active_thread[(101*4)+2] <= 1'b0;
                  active_thread[(101*4)+3] <= 1'b0;
                  spc101_inst_done         <= 0;
                  spc101_phy_pc_w          <= 0;
                end else begin
                  active_thread[(101*4)]   <= 1'b1;
                  active_thread[(101*4)+1] <= 1'b1;
                  active_thread[(101*4)+2] <= 1'b1;
                  active_thread[(101*4)+3] <= 1'b1;
                  spc101_inst_done         <= `ARIANE_CORE101.piton_pc_vld;
                  spc101_phy_pc_w          <= `ARIANE_CORE101.piton_pc;
                end
            end
    

            assign spc102_thread_id = 2'b00;
            assign spc102_rtl_pc = spc102_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(102*4)]   <= 1'b0;
                  active_thread[(102*4)+1] <= 1'b0;
                  active_thread[(102*4)+2] <= 1'b0;
                  active_thread[(102*4)+3] <= 1'b0;
                  spc102_inst_done         <= 0;
                  spc102_phy_pc_w          <= 0;
                end else begin
                  active_thread[(102*4)]   <= 1'b1;
                  active_thread[(102*4)+1] <= 1'b1;
                  active_thread[(102*4)+2] <= 1'b1;
                  active_thread[(102*4)+3] <= 1'b1;
                  spc102_inst_done         <= `ARIANE_CORE102.piton_pc_vld;
                  spc102_phy_pc_w          <= `ARIANE_CORE102.piton_pc;
                end
            end
    

            assign spc103_thread_id = 2'b00;
            assign spc103_rtl_pc = spc103_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(103*4)]   <= 1'b0;
                  active_thread[(103*4)+1] <= 1'b0;
                  active_thread[(103*4)+2] <= 1'b0;
                  active_thread[(103*4)+3] <= 1'b0;
                  spc103_inst_done         <= 0;
                  spc103_phy_pc_w          <= 0;
                end else begin
                  active_thread[(103*4)]   <= 1'b1;
                  active_thread[(103*4)+1] <= 1'b1;
                  active_thread[(103*4)+2] <= 1'b1;
                  active_thread[(103*4)+3] <= 1'b1;
                  spc103_inst_done         <= `ARIANE_CORE103.piton_pc_vld;
                  spc103_phy_pc_w          <= `ARIANE_CORE103.piton_pc;
                end
            end
    

            assign spc104_thread_id = 2'b00;
            assign spc104_rtl_pc = spc104_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(104*4)]   <= 1'b0;
                  active_thread[(104*4)+1] <= 1'b0;
                  active_thread[(104*4)+2] <= 1'b0;
                  active_thread[(104*4)+3] <= 1'b0;
                  spc104_inst_done         <= 0;
                  spc104_phy_pc_w          <= 0;
                end else begin
                  active_thread[(104*4)]   <= 1'b1;
                  active_thread[(104*4)+1] <= 1'b1;
                  active_thread[(104*4)+2] <= 1'b1;
                  active_thread[(104*4)+3] <= 1'b1;
                  spc104_inst_done         <= `ARIANE_CORE104.piton_pc_vld;
                  spc104_phy_pc_w          <= `ARIANE_CORE104.piton_pc;
                end
            end
    

            assign spc105_thread_id = 2'b00;
            assign spc105_rtl_pc = spc105_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(105*4)]   <= 1'b0;
                  active_thread[(105*4)+1] <= 1'b0;
                  active_thread[(105*4)+2] <= 1'b0;
                  active_thread[(105*4)+3] <= 1'b0;
                  spc105_inst_done         <= 0;
                  spc105_phy_pc_w          <= 0;
                end else begin
                  active_thread[(105*4)]   <= 1'b1;
                  active_thread[(105*4)+1] <= 1'b1;
                  active_thread[(105*4)+2] <= 1'b1;
                  active_thread[(105*4)+3] <= 1'b1;
                  spc105_inst_done         <= `ARIANE_CORE105.piton_pc_vld;
                  spc105_phy_pc_w          <= `ARIANE_CORE105.piton_pc;
                end
            end
    

            assign spc106_thread_id = 2'b00;
            assign spc106_rtl_pc = spc106_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(106*4)]   <= 1'b0;
                  active_thread[(106*4)+1] <= 1'b0;
                  active_thread[(106*4)+2] <= 1'b0;
                  active_thread[(106*4)+3] <= 1'b0;
                  spc106_inst_done         <= 0;
                  spc106_phy_pc_w          <= 0;
                end else begin
                  active_thread[(106*4)]   <= 1'b1;
                  active_thread[(106*4)+1] <= 1'b1;
                  active_thread[(106*4)+2] <= 1'b1;
                  active_thread[(106*4)+3] <= 1'b1;
                  spc106_inst_done         <= `ARIANE_CORE106.piton_pc_vld;
                  spc106_phy_pc_w          <= `ARIANE_CORE106.piton_pc;
                end
            end
    

            assign spc107_thread_id = 2'b00;
            assign spc107_rtl_pc = spc107_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(107*4)]   <= 1'b0;
                  active_thread[(107*4)+1] <= 1'b0;
                  active_thread[(107*4)+2] <= 1'b0;
                  active_thread[(107*4)+3] <= 1'b0;
                  spc107_inst_done         <= 0;
                  spc107_phy_pc_w          <= 0;
                end else begin
                  active_thread[(107*4)]   <= 1'b1;
                  active_thread[(107*4)+1] <= 1'b1;
                  active_thread[(107*4)+2] <= 1'b1;
                  active_thread[(107*4)+3] <= 1'b1;
                  spc107_inst_done         <= `ARIANE_CORE107.piton_pc_vld;
                  spc107_phy_pc_w          <= `ARIANE_CORE107.piton_pc;
                end
            end
    

            assign spc108_thread_id = 2'b00;
            assign spc108_rtl_pc = spc108_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(108*4)]   <= 1'b0;
                  active_thread[(108*4)+1] <= 1'b0;
                  active_thread[(108*4)+2] <= 1'b0;
                  active_thread[(108*4)+3] <= 1'b0;
                  spc108_inst_done         <= 0;
                  spc108_phy_pc_w          <= 0;
                end else begin
                  active_thread[(108*4)]   <= 1'b1;
                  active_thread[(108*4)+1] <= 1'b1;
                  active_thread[(108*4)+2] <= 1'b1;
                  active_thread[(108*4)+3] <= 1'b1;
                  spc108_inst_done         <= `ARIANE_CORE108.piton_pc_vld;
                  spc108_phy_pc_w          <= `ARIANE_CORE108.piton_pc;
                end
            end
    

            assign spc109_thread_id = 2'b00;
            assign spc109_rtl_pc = spc109_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(109*4)]   <= 1'b0;
                  active_thread[(109*4)+1] <= 1'b0;
                  active_thread[(109*4)+2] <= 1'b0;
                  active_thread[(109*4)+3] <= 1'b0;
                  spc109_inst_done         <= 0;
                  spc109_phy_pc_w          <= 0;
                end else begin
                  active_thread[(109*4)]   <= 1'b1;
                  active_thread[(109*4)+1] <= 1'b1;
                  active_thread[(109*4)+2] <= 1'b1;
                  active_thread[(109*4)+3] <= 1'b1;
                  spc109_inst_done         <= `ARIANE_CORE109.piton_pc_vld;
                  spc109_phy_pc_w          <= `ARIANE_CORE109.piton_pc;
                end
            end
    

            assign spc110_thread_id = 2'b00;
            assign spc110_rtl_pc = spc110_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(110*4)]   <= 1'b0;
                  active_thread[(110*4)+1] <= 1'b0;
                  active_thread[(110*4)+2] <= 1'b0;
                  active_thread[(110*4)+3] <= 1'b0;
                  spc110_inst_done         <= 0;
                  spc110_phy_pc_w          <= 0;
                end else begin
                  active_thread[(110*4)]   <= 1'b1;
                  active_thread[(110*4)+1] <= 1'b1;
                  active_thread[(110*4)+2] <= 1'b1;
                  active_thread[(110*4)+3] <= 1'b1;
                  spc110_inst_done         <= `ARIANE_CORE110.piton_pc_vld;
                  spc110_phy_pc_w          <= `ARIANE_CORE110.piton_pc;
                end
            end
    

            assign spc111_thread_id = 2'b00;
            assign spc111_rtl_pc = spc111_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(111*4)]   <= 1'b0;
                  active_thread[(111*4)+1] <= 1'b0;
                  active_thread[(111*4)+2] <= 1'b0;
                  active_thread[(111*4)+3] <= 1'b0;
                  spc111_inst_done         <= 0;
                  spc111_phy_pc_w          <= 0;
                end else begin
                  active_thread[(111*4)]   <= 1'b1;
                  active_thread[(111*4)+1] <= 1'b1;
                  active_thread[(111*4)+2] <= 1'b1;
                  active_thread[(111*4)+3] <= 1'b1;
                  spc111_inst_done         <= `ARIANE_CORE111.piton_pc_vld;
                  spc111_phy_pc_w          <= `ARIANE_CORE111.piton_pc;
                end
            end
    

            assign spc112_thread_id = 2'b00;
            assign spc112_rtl_pc = spc112_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(112*4)]   <= 1'b0;
                  active_thread[(112*4)+1] <= 1'b0;
                  active_thread[(112*4)+2] <= 1'b0;
                  active_thread[(112*4)+3] <= 1'b0;
                  spc112_inst_done         <= 0;
                  spc112_phy_pc_w          <= 0;
                end else begin
                  active_thread[(112*4)]   <= 1'b1;
                  active_thread[(112*4)+1] <= 1'b1;
                  active_thread[(112*4)+2] <= 1'b1;
                  active_thread[(112*4)+3] <= 1'b1;
                  spc112_inst_done         <= `ARIANE_CORE112.piton_pc_vld;
                  spc112_phy_pc_w          <= `ARIANE_CORE112.piton_pc;
                end
            end
    

            assign spc113_thread_id = 2'b00;
            assign spc113_rtl_pc = spc113_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(113*4)]   <= 1'b0;
                  active_thread[(113*4)+1] <= 1'b0;
                  active_thread[(113*4)+2] <= 1'b0;
                  active_thread[(113*4)+3] <= 1'b0;
                  spc113_inst_done         <= 0;
                  spc113_phy_pc_w          <= 0;
                end else begin
                  active_thread[(113*4)]   <= 1'b1;
                  active_thread[(113*4)+1] <= 1'b1;
                  active_thread[(113*4)+2] <= 1'b1;
                  active_thread[(113*4)+3] <= 1'b1;
                  spc113_inst_done         <= `ARIANE_CORE113.piton_pc_vld;
                  spc113_phy_pc_w          <= `ARIANE_CORE113.piton_pc;
                end
            end
    

            assign spc114_thread_id = 2'b00;
            assign spc114_rtl_pc = spc114_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(114*4)]   <= 1'b0;
                  active_thread[(114*4)+1] <= 1'b0;
                  active_thread[(114*4)+2] <= 1'b0;
                  active_thread[(114*4)+3] <= 1'b0;
                  spc114_inst_done         <= 0;
                  spc114_phy_pc_w          <= 0;
                end else begin
                  active_thread[(114*4)]   <= 1'b1;
                  active_thread[(114*4)+1] <= 1'b1;
                  active_thread[(114*4)+2] <= 1'b1;
                  active_thread[(114*4)+3] <= 1'b1;
                  spc114_inst_done         <= `ARIANE_CORE114.piton_pc_vld;
                  spc114_phy_pc_w          <= `ARIANE_CORE114.piton_pc;
                end
            end
    

            assign spc115_thread_id = 2'b00;
            assign spc115_rtl_pc = spc115_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(115*4)]   <= 1'b0;
                  active_thread[(115*4)+1] <= 1'b0;
                  active_thread[(115*4)+2] <= 1'b0;
                  active_thread[(115*4)+3] <= 1'b0;
                  spc115_inst_done         <= 0;
                  spc115_phy_pc_w          <= 0;
                end else begin
                  active_thread[(115*4)]   <= 1'b1;
                  active_thread[(115*4)+1] <= 1'b1;
                  active_thread[(115*4)+2] <= 1'b1;
                  active_thread[(115*4)+3] <= 1'b1;
                  spc115_inst_done         <= `ARIANE_CORE115.piton_pc_vld;
                  spc115_phy_pc_w          <= `ARIANE_CORE115.piton_pc;
                end
            end
    

            assign spc116_thread_id = 2'b00;
            assign spc116_rtl_pc = spc116_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(116*4)]   <= 1'b0;
                  active_thread[(116*4)+1] <= 1'b0;
                  active_thread[(116*4)+2] <= 1'b0;
                  active_thread[(116*4)+3] <= 1'b0;
                  spc116_inst_done         <= 0;
                  spc116_phy_pc_w          <= 0;
                end else begin
                  active_thread[(116*4)]   <= 1'b1;
                  active_thread[(116*4)+1] <= 1'b1;
                  active_thread[(116*4)+2] <= 1'b1;
                  active_thread[(116*4)+3] <= 1'b1;
                  spc116_inst_done         <= `ARIANE_CORE116.piton_pc_vld;
                  spc116_phy_pc_w          <= `ARIANE_CORE116.piton_pc;
                end
            end
    

            assign spc117_thread_id = 2'b00;
            assign spc117_rtl_pc = spc117_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(117*4)]   <= 1'b0;
                  active_thread[(117*4)+1] <= 1'b0;
                  active_thread[(117*4)+2] <= 1'b0;
                  active_thread[(117*4)+3] <= 1'b0;
                  spc117_inst_done         <= 0;
                  spc117_phy_pc_w          <= 0;
                end else begin
                  active_thread[(117*4)]   <= 1'b1;
                  active_thread[(117*4)+1] <= 1'b1;
                  active_thread[(117*4)+2] <= 1'b1;
                  active_thread[(117*4)+3] <= 1'b1;
                  spc117_inst_done         <= `ARIANE_CORE117.piton_pc_vld;
                  spc117_phy_pc_w          <= `ARIANE_CORE117.piton_pc;
                end
            end
    

            assign spc118_thread_id = 2'b00;
            assign spc118_rtl_pc = spc118_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(118*4)]   <= 1'b0;
                  active_thread[(118*4)+1] <= 1'b0;
                  active_thread[(118*4)+2] <= 1'b0;
                  active_thread[(118*4)+3] <= 1'b0;
                  spc118_inst_done         <= 0;
                  spc118_phy_pc_w          <= 0;
                end else begin
                  active_thread[(118*4)]   <= 1'b1;
                  active_thread[(118*4)+1] <= 1'b1;
                  active_thread[(118*4)+2] <= 1'b1;
                  active_thread[(118*4)+3] <= 1'b1;
                  spc118_inst_done         <= `ARIANE_CORE118.piton_pc_vld;
                  spc118_phy_pc_w          <= `ARIANE_CORE118.piton_pc;
                end
            end
    

            assign spc119_thread_id = 2'b00;
            assign spc119_rtl_pc = spc119_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(119*4)]   <= 1'b0;
                  active_thread[(119*4)+1] <= 1'b0;
                  active_thread[(119*4)+2] <= 1'b0;
                  active_thread[(119*4)+3] <= 1'b0;
                  spc119_inst_done         <= 0;
                  spc119_phy_pc_w          <= 0;
                end else begin
                  active_thread[(119*4)]   <= 1'b1;
                  active_thread[(119*4)+1] <= 1'b1;
                  active_thread[(119*4)+2] <= 1'b1;
                  active_thread[(119*4)+3] <= 1'b1;
                  spc119_inst_done         <= `ARIANE_CORE119.piton_pc_vld;
                  spc119_phy_pc_w          <= `ARIANE_CORE119.piton_pc;
                end
            end
    

            assign spc120_thread_id = 2'b00;
            assign spc120_rtl_pc = spc120_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(120*4)]   <= 1'b0;
                  active_thread[(120*4)+1] <= 1'b0;
                  active_thread[(120*4)+2] <= 1'b0;
                  active_thread[(120*4)+3] <= 1'b0;
                  spc120_inst_done         <= 0;
                  spc120_phy_pc_w          <= 0;
                end else begin
                  active_thread[(120*4)]   <= 1'b1;
                  active_thread[(120*4)+1] <= 1'b1;
                  active_thread[(120*4)+2] <= 1'b1;
                  active_thread[(120*4)+3] <= 1'b1;
                  spc120_inst_done         <= `ARIANE_CORE120.piton_pc_vld;
                  spc120_phy_pc_w          <= `ARIANE_CORE120.piton_pc;
                end
            end
    

            assign spc121_thread_id = 2'b00;
            assign spc121_rtl_pc = spc121_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(121*4)]   <= 1'b0;
                  active_thread[(121*4)+1] <= 1'b0;
                  active_thread[(121*4)+2] <= 1'b0;
                  active_thread[(121*4)+3] <= 1'b0;
                  spc121_inst_done         <= 0;
                  spc121_phy_pc_w          <= 0;
                end else begin
                  active_thread[(121*4)]   <= 1'b1;
                  active_thread[(121*4)+1] <= 1'b1;
                  active_thread[(121*4)+2] <= 1'b1;
                  active_thread[(121*4)+3] <= 1'b1;
                  spc121_inst_done         <= `ARIANE_CORE121.piton_pc_vld;
                  spc121_phy_pc_w          <= `ARIANE_CORE121.piton_pc;
                end
            end
    

            assign spc122_thread_id = 2'b00;
            assign spc122_rtl_pc = spc122_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(122*4)]   <= 1'b0;
                  active_thread[(122*4)+1] <= 1'b0;
                  active_thread[(122*4)+2] <= 1'b0;
                  active_thread[(122*4)+3] <= 1'b0;
                  spc122_inst_done         <= 0;
                  spc122_phy_pc_w          <= 0;
                end else begin
                  active_thread[(122*4)]   <= 1'b1;
                  active_thread[(122*4)+1] <= 1'b1;
                  active_thread[(122*4)+2] <= 1'b1;
                  active_thread[(122*4)+3] <= 1'b1;
                  spc122_inst_done         <= `ARIANE_CORE122.piton_pc_vld;
                  spc122_phy_pc_w          <= `ARIANE_CORE122.piton_pc;
                end
            end
    

            assign spc123_thread_id = 2'b00;
            assign spc123_rtl_pc = spc123_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(123*4)]   <= 1'b0;
                  active_thread[(123*4)+1] <= 1'b0;
                  active_thread[(123*4)+2] <= 1'b0;
                  active_thread[(123*4)+3] <= 1'b0;
                  spc123_inst_done         <= 0;
                  spc123_phy_pc_w          <= 0;
                end else begin
                  active_thread[(123*4)]   <= 1'b1;
                  active_thread[(123*4)+1] <= 1'b1;
                  active_thread[(123*4)+2] <= 1'b1;
                  active_thread[(123*4)+3] <= 1'b1;
                  spc123_inst_done         <= `ARIANE_CORE123.piton_pc_vld;
                  spc123_phy_pc_w          <= `ARIANE_CORE123.piton_pc;
                end
            end
    

            assign spc124_thread_id = 2'b00;
            assign spc124_rtl_pc = spc124_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(124*4)]   <= 1'b0;
                  active_thread[(124*4)+1] <= 1'b0;
                  active_thread[(124*4)+2] <= 1'b0;
                  active_thread[(124*4)+3] <= 1'b0;
                  spc124_inst_done         <= 0;
                  spc124_phy_pc_w          <= 0;
                end else begin
                  active_thread[(124*4)]   <= 1'b1;
                  active_thread[(124*4)+1] <= 1'b1;
                  active_thread[(124*4)+2] <= 1'b1;
                  active_thread[(124*4)+3] <= 1'b1;
                  spc124_inst_done         <= `ARIANE_CORE124.piton_pc_vld;
                  spc124_phy_pc_w          <= `ARIANE_CORE124.piton_pc;
                end
            end
    

            assign spc125_thread_id = 2'b00;
            assign spc125_rtl_pc = spc125_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(125*4)]   <= 1'b0;
                  active_thread[(125*4)+1] <= 1'b0;
                  active_thread[(125*4)+2] <= 1'b0;
                  active_thread[(125*4)+3] <= 1'b0;
                  spc125_inst_done         <= 0;
                  spc125_phy_pc_w          <= 0;
                end else begin
                  active_thread[(125*4)]   <= 1'b1;
                  active_thread[(125*4)+1] <= 1'b1;
                  active_thread[(125*4)+2] <= 1'b1;
                  active_thread[(125*4)+3] <= 1'b1;
                  spc125_inst_done         <= `ARIANE_CORE125.piton_pc_vld;
                  spc125_phy_pc_w          <= `ARIANE_CORE125.piton_pc;
                end
            end
    

            assign spc126_thread_id = 2'b00;
            assign spc126_rtl_pc = spc126_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(126*4)]   <= 1'b0;
                  active_thread[(126*4)+1] <= 1'b0;
                  active_thread[(126*4)+2] <= 1'b0;
                  active_thread[(126*4)+3] <= 1'b0;
                  spc126_inst_done         <= 0;
                  spc126_phy_pc_w          <= 0;
                end else begin
                  active_thread[(126*4)]   <= 1'b1;
                  active_thread[(126*4)+1] <= 1'b1;
                  active_thread[(126*4)+2] <= 1'b1;
                  active_thread[(126*4)+3] <= 1'b1;
                  spc126_inst_done         <= `ARIANE_CORE126.piton_pc_vld;
                  spc126_phy_pc_w          <= `ARIANE_CORE126.piton_pc;
                end
            end
    

            assign spc127_thread_id = 2'b00;
            assign spc127_rtl_pc = spc127_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(127*4)]   <= 1'b0;
                  active_thread[(127*4)+1] <= 1'b0;
                  active_thread[(127*4)+2] <= 1'b0;
                  active_thread[(127*4)+3] <= 1'b0;
                  spc127_inst_done         <= 0;
                  spc127_phy_pc_w          <= 0;
                end else begin
                  active_thread[(127*4)]   <= 1'b1;
                  active_thread[(127*4)+1] <= 1'b1;
                  active_thread[(127*4)+2] <= 1'b1;
                  active_thread[(127*4)+3] <= 1'b1;
                  spc127_inst_done         <= `ARIANE_CORE127.piton_pc_vld;
                  spc127_phy_pc_w          <= `ARIANE_CORE127.piton_pc;
                end
            end
    

            assign spc128_thread_id = 2'b00;
            assign spc128_rtl_pc = spc128_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(128*4)]   <= 1'b0;
                  active_thread[(128*4)+1] <= 1'b0;
                  active_thread[(128*4)+2] <= 1'b0;
                  active_thread[(128*4)+3] <= 1'b0;
                  spc128_inst_done         <= 0;
                  spc128_phy_pc_w          <= 0;
                end else begin
                  active_thread[(128*4)]   <= 1'b1;
                  active_thread[(128*4)+1] <= 1'b1;
                  active_thread[(128*4)+2] <= 1'b1;
                  active_thread[(128*4)+3] <= 1'b1;
                  spc128_inst_done         <= `ARIANE_CORE128.piton_pc_vld;
                  spc128_phy_pc_w          <= `ARIANE_CORE128.piton_pc;
                end
            end
    

            assign spc129_thread_id = 2'b00;
            assign spc129_rtl_pc = spc129_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(129*4)]   <= 1'b0;
                  active_thread[(129*4)+1] <= 1'b0;
                  active_thread[(129*4)+2] <= 1'b0;
                  active_thread[(129*4)+3] <= 1'b0;
                  spc129_inst_done         <= 0;
                  spc129_phy_pc_w          <= 0;
                end else begin
                  active_thread[(129*4)]   <= 1'b1;
                  active_thread[(129*4)+1] <= 1'b1;
                  active_thread[(129*4)+2] <= 1'b1;
                  active_thread[(129*4)+3] <= 1'b1;
                  spc129_inst_done         <= `ARIANE_CORE129.piton_pc_vld;
                  spc129_phy_pc_w          <= `ARIANE_CORE129.piton_pc;
                end
            end
    

            assign spc130_thread_id = 2'b00;
            assign spc130_rtl_pc = spc130_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(130*4)]   <= 1'b0;
                  active_thread[(130*4)+1] <= 1'b0;
                  active_thread[(130*4)+2] <= 1'b0;
                  active_thread[(130*4)+3] <= 1'b0;
                  spc130_inst_done         <= 0;
                  spc130_phy_pc_w          <= 0;
                end else begin
                  active_thread[(130*4)]   <= 1'b1;
                  active_thread[(130*4)+1] <= 1'b1;
                  active_thread[(130*4)+2] <= 1'b1;
                  active_thread[(130*4)+3] <= 1'b1;
                  spc130_inst_done         <= `ARIANE_CORE130.piton_pc_vld;
                  spc130_phy_pc_w          <= `ARIANE_CORE130.piton_pc;
                end
            end
    

            assign spc131_thread_id = 2'b00;
            assign spc131_rtl_pc = spc131_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(131*4)]   <= 1'b0;
                  active_thread[(131*4)+1] <= 1'b0;
                  active_thread[(131*4)+2] <= 1'b0;
                  active_thread[(131*4)+3] <= 1'b0;
                  spc131_inst_done         <= 0;
                  spc131_phy_pc_w          <= 0;
                end else begin
                  active_thread[(131*4)]   <= 1'b1;
                  active_thread[(131*4)+1] <= 1'b1;
                  active_thread[(131*4)+2] <= 1'b1;
                  active_thread[(131*4)+3] <= 1'b1;
                  spc131_inst_done         <= `ARIANE_CORE131.piton_pc_vld;
                  spc131_phy_pc_w          <= `ARIANE_CORE131.piton_pc;
                end
            end
    

            assign spc132_thread_id = 2'b00;
            assign spc132_rtl_pc = spc132_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(132*4)]   <= 1'b0;
                  active_thread[(132*4)+1] <= 1'b0;
                  active_thread[(132*4)+2] <= 1'b0;
                  active_thread[(132*4)+3] <= 1'b0;
                  spc132_inst_done         <= 0;
                  spc132_phy_pc_w          <= 0;
                end else begin
                  active_thread[(132*4)]   <= 1'b1;
                  active_thread[(132*4)+1] <= 1'b1;
                  active_thread[(132*4)+2] <= 1'b1;
                  active_thread[(132*4)+3] <= 1'b1;
                  spc132_inst_done         <= `ARIANE_CORE132.piton_pc_vld;
                  spc132_phy_pc_w          <= `ARIANE_CORE132.piton_pc;
                end
            end
    

            assign spc133_thread_id = 2'b00;
            assign spc133_rtl_pc = spc133_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(133*4)]   <= 1'b0;
                  active_thread[(133*4)+1] <= 1'b0;
                  active_thread[(133*4)+2] <= 1'b0;
                  active_thread[(133*4)+3] <= 1'b0;
                  spc133_inst_done         <= 0;
                  spc133_phy_pc_w          <= 0;
                end else begin
                  active_thread[(133*4)]   <= 1'b1;
                  active_thread[(133*4)+1] <= 1'b1;
                  active_thread[(133*4)+2] <= 1'b1;
                  active_thread[(133*4)+3] <= 1'b1;
                  spc133_inst_done         <= `ARIANE_CORE133.piton_pc_vld;
                  spc133_phy_pc_w          <= `ARIANE_CORE133.piton_pc;
                end
            end
    

            assign spc134_thread_id = 2'b00;
            assign spc134_rtl_pc = spc134_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(134*4)]   <= 1'b0;
                  active_thread[(134*4)+1] <= 1'b0;
                  active_thread[(134*4)+2] <= 1'b0;
                  active_thread[(134*4)+3] <= 1'b0;
                  spc134_inst_done         <= 0;
                  spc134_phy_pc_w          <= 0;
                end else begin
                  active_thread[(134*4)]   <= 1'b1;
                  active_thread[(134*4)+1] <= 1'b1;
                  active_thread[(134*4)+2] <= 1'b1;
                  active_thread[(134*4)+3] <= 1'b1;
                  spc134_inst_done         <= `ARIANE_CORE134.piton_pc_vld;
                  spc134_phy_pc_w          <= `ARIANE_CORE134.piton_pc;
                end
            end
    

            assign spc135_thread_id = 2'b00;
            assign spc135_rtl_pc = spc135_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(135*4)]   <= 1'b0;
                  active_thread[(135*4)+1] <= 1'b0;
                  active_thread[(135*4)+2] <= 1'b0;
                  active_thread[(135*4)+3] <= 1'b0;
                  spc135_inst_done         <= 0;
                  spc135_phy_pc_w          <= 0;
                end else begin
                  active_thread[(135*4)]   <= 1'b1;
                  active_thread[(135*4)+1] <= 1'b1;
                  active_thread[(135*4)+2] <= 1'b1;
                  active_thread[(135*4)+3] <= 1'b1;
                  spc135_inst_done         <= `ARIANE_CORE135.piton_pc_vld;
                  spc135_phy_pc_w          <= `ARIANE_CORE135.piton_pc;
                end
            end
    

            assign spc136_thread_id = 2'b00;
            assign spc136_rtl_pc = spc136_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(136*4)]   <= 1'b0;
                  active_thread[(136*4)+1] <= 1'b0;
                  active_thread[(136*4)+2] <= 1'b0;
                  active_thread[(136*4)+3] <= 1'b0;
                  spc136_inst_done         <= 0;
                  spc136_phy_pc_w          <= 0;
                end else begin
                  active_thread[(136*4)]   <= 1'b1;
                  active_thread[(136*4)+1] <= 1'b1;
                  active_thread[(136*4)+2] <= 1'b1;
                  active_thread[(136*4)+3] <= 1'b1;
                  spc136_inst_done         <= `ARIANE_CORE136.piton_pc_vld;
                  spc136_phy_pc_w          <= `ARIANE_CORE136.piton_pc;
                end
            end
    

            assign spc137_thread_id = 2'b00;
            assign spc137_rtl_pc = spc137_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(137*4)]   <= 1'b0;
                  active_thread[(137*4)+1] <= 1'b0;
                  active_thread[(137*4)+2] <= 1'b0;
                  active_thread[(137*4)+3] <= 1'b0;
                  spc137_inst_done         <= 0;
                  spc137_phy_pc_w          <= 0;
                end else begin
                  active_thread[(137*4)]   <= 1'b1;
                  active_thread[(137*4)+1] <= 1'b1;
                  active_thread[(137*4)+2] <= 1'b1;
                  active_thread[(137*4)+3] <= 1'b1;
                  spc137_inst_done         <= `ARIANE_CORE137.piton_pc_vld;
                  spc137_phy_pc_w          <= `ARIANE_CORE137.piton_pc;
                end
            end
    

            assign spc138_thread_id = 2'b00;
            assign spc138_rtl_pc = spc138_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(138*4)]   <= 1'b0;
                  active_thread[(138*4)+1] <= 1'b0;
                  active_thread[(138*4)+2] <= 1'b0;
                  active_thread[(138*4)+3] <= 1'b0;
                  spc138_inst_done         <= 0;
                  spc138_phy_pc_w          <= 0;
                end else begin
                  active_thread[(138*4)]   <= 1'b1;
                  active_thread[(138*4)+1] <= 1'b1;
                  active_thread[(138*4)+2] <= 1'b1;
                  active_thread[(138*4)+3] <= 1'b1;
                  spc138_inst_done         <= `ARIANE_CORE138.piton_pc_vld;
                  spc138_phy_pc_w          <= `ARIANE_CORE138.piton_pc;
                end
            end
    

            assign spc139_thread_id = 2'b00;
            assign spc139_rtl_pc = spc139_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(139*4)]   <= 1'b0;
                  active_thread[(139*4)+1] <= 1'b0;
                  active_thread[(139*4)+2] <= 1'b0;
                  active_thread[(139*4)+3] <= 1'b0;
                  spc139_inst_done         <= 0;
                  spc139_phy_pc_w          <= 0;
                end else begin
                  active_thread[(139*4)]   <= 1'b1;
                  active_thread[(139*4)+1] <= 1'b1;
                  active_thread[(139*4)+2] <= 1'b1;
                  active_thread[(139*4)+3] <= 1'b1;
                  spc139_inst_done         <= `ARIANE_CORE139.piton_pc_vld;
                  spc139_phy_pc_w          <= `ARIANE_CORE139.piton_pc;
                end
            end
    

            assign spc140_thread_id = 2'b00;
            assign spc140_rtl_pc = spc140_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(140*4)]   <= 1'b0;
                  active_thread[(140*4)+1] <= 1'b0;
                  active_thread[(140*4)+2] <= 1'b0;
                  active_thread[(140*4)+3] <= 1'b0;
                  spc140_inst_done         <= 0;
                  spc140_phy_pc_w          <= 0;
                end else begin
                  active_thread[(140*4)]   <= 1'b1;
                  active_thread[(140*4)+1] <= 1'b1;
                  active_thread[(140*4)+2] <= 1'b1;
                  active_thread[(140*4)+3] <= 1'b1;
                  spc140_inst_done         <= `ARIANE_CORE140.piton_pc_vld;
                  spc140_phy_pc_w          <= `ARIANE_CORE140.piton_pc;
                end
            end
    

            assign spc141_thread_id = 2'b00;
            assign spc141_rtl_pc = spc141_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(141*4)]   <= 1'b0;
                  active_thread[(141*4)+1] <= 1'b0;
                  active_thread[(141*4)+2] <= 1'b0;
                  active_thread[(141*4)+3] <= 1'b0;
                  spc141_inst_done         <= 0;
                  spc141_phy_pc_w          <= 0;
                end else begin
                  active_thread[(141*4)]   <= 1'b1;
                  active_thread[(141*4)+1] <= 1'b1;
                  active_thread[(141*4)+2] <= 1'b1;
                  active_thread[(141*4)+3] <= 1'b1;
                  spc141_inst_done         <= `ARIANE_CORE141.piton_pc_vld;
                  spc141_phy_pc_w          <= `ARIANE_CORE141.piton_pc;
                end
            end
    

            assign spc142_thread_id = 2'b00;
            assign spc142_rtl_pc = spc142_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(142*4)]   <= 1'b0;
                  active_thread[(142*4)+1] <= 1'b0;
                  active_thread[(142*4)+2] <= 1'b0;
                  active_thread[(142*4)+3] <= 1'b0;
                  spc142_inst_done         <= 0;
                  spc142_phy_pc_w          <= 0;
                end else begin
                  active_thread[(142*4)]   <= 1'b1;
                  active_thread[(142*4)+1] <= 1'b1;
                  active_thread[(142*4)+2] <= 1'b1;
                  active_thread[(142*4)+3] <= 1'b1;
                  spc142_inst_done         <= `ARIANE_CORE142.piton_pc_vld;
                  spc142_phy_pc_w          <= `ARIANE_CORE142.piton_pc;
                end
            end
    

            assign spc143_thread_id = 2'b00;
            assign spc143_rtl_pc = spc143_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(143*4)]   <= 1'b0;
                  active_thread[(143*4)+1] <= 1'b0;
                  active_thread[(143*4)+2] <= 1'b0;
                  active_thread[(143*4)+3] <= 1'b0;
                  spc143_inst_done         <= 0;
                  spc143_phy_pc_w          <= 0;
                end else begin
                  active_thread[(143*4)]   <= 1'b1;
                  active_thread[(143*4)+1] <= 1'b1;
                  active_thread[(143*4)+2] <= 1'b1;
                  active_thread[(143*4)+3] <= 1'b1;
                  spc143_inst_done         <= `ARIANE_CORE143.piton_pc_vld;
                  spc143_phy_pc_w          <= `ARIANE_CORE143.piton_pc;
                end
            end
    

            assign spc144_thread_id = 2'b00;
            assign spc144_rtl_pc = spc144_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(144*4)]   <= 1'b0;
                  active_thread[(144*4)+1] <= 1'b0;
                  active_thread[(144*4)+2] <= 1'b0;
                  active_thread[(144*4)+3] <= 1'b0;
                  spc144_inst_done         <= 0;
                  spc144_phy_pc_w          <= 0;
                end else begin
                  active_thread[(144*4)]   <= 1'b1;
                  active_thread[(144*4)+1] <= 1'b1;
                  active_thread[(144*4)+2] <= 1'b1;
                  active_thread[(144*4)+3] <= 1'b1;
                  spc144_inst_done         <= `ARIANE_CORE144.piton_pc_vld;
                  spc144_phy_pc_w          <= `ARIANE_CORE144.piton_pc;
                end
            end
    

            assign spc145_thread_id = 2'b00;
            assign spc145_rtl_pc = spc145_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(145*4)]   <= 1'b0;
                  active_thread[(145*4)+1] <= 1'b0;
                  active_thread[(145*4)+2] <= 1'b0;
                  active_thread[(145*4)+3] <= 1'b0;
                  spc145_inst_done         <= 0;
                  spc145_phy_pc_w          <= 0;
                end else begin
                  active_thread[(145*4)]   <= 1'b1;
                  active_thread[(145*4)+1] <= 1'b1;
                  active_thread[(145*4)+2] <= 1'b1;
                  active_thread[(145*4)+3] <= 1'b1;
                  spc145_inst_done         <= `ARIANE_CORE145.piton_pc_vld;
                  spc145_phy_pc_w          <= `ARIANE_CORE145.piton_pc;
                end
            end
    

            assign spc146_thread_id = 2'b00;
            assign spc146_rtl_pc = spc146_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(146*4)]   <= 1'b0;
                  active_thread[(146*4)+1] <= 1'b0;
                  active_thread[(146*4)+2] <= 1'b0;
                  active_thread[(146*4)+3] <= 1'b0;
                  spc146_inst_done         <= 0;
                  spc146_phy_pc_w          <= 0;
                end else begin
                  active_thread[(146*4)]   <= 1'b1;
                  active_thread[(146*4)+1] <= 1'b1;
                  active_thread[(146*4)+2] <= 1'b1;
                  active_thread[(146*4)+3] <= 1'b1;
                  spc146_inst_done         <= `ARIANE_CORE146.piton_pc_vld;
                  spc146_phy_pc_w          <= `ARIANE_CORE146.piton_pc;
                end
            end
    

            assign spc147_thread_id = 2'b00;
            assign spc147_rtl_pc = spc147_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(147*4)]   <= 1'b0;
                  active_thread[(147*4)+1] <= 1'b0;
                  active_thread[(147*4)+2] <= 1'b0;
                  active_thread[(147*4)+3] <= 1'b0;
                  spc147_inst_done         <= 0;
                  spc147_phy_pc_w          <= 0;
                end else begin
                  active_thread[(147*4)]   <= 1'b1;
                  active_thread[(147*4)+1] <= 1'b1;
                  active_thread[(147*4)+2] <= 1'b1;
                  active_thread[(147*4)+3] <= 1'b1;
                  spc147_inst_done         <= `ARIANE_CORE147.piton_pc_vld;
                  spc147_phy_pc_w          <= `ARIANE_CORE147.piton_pc;
                end
            end
    

            assign spc148_thread_id = 2'b00;
            assign spc148_rtl_pc = spc148_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(148*4)]   <= 1'b0;
                  active_thread[(148*4)+1] <= 1'b0;
                  active_thread[(148*4)+2] <= 1'b0;
                  active_thread[(148*4)+3] <= 1'b0;
                  spc148_inst_done         <= 0;
                  spc148_phy_pc_w          <= 0;
                end else begin
                  active_thread[(148*4)]   <= 1'b1;
                  active_thread[(148*4)+1] <= 1'b1;
                  active_thread[(148*4)+2] <= 1'b1;
                  active_thread[(148*4)+3] <= 1'b1;
                  spc148_inst_done         <= `ARIANE_CORE148.piton_pc_vld;
                  spc148_phy_pc_w          <= `ARIANE_CORE148.piton_pc;
                end
            end
    

            assign spc149_thread_id = 2'b00;
            assign spc149_rtl_pc = spc149_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(149*4)]   <= 1'b0;
                  active_thread[(149*4)+1] <= 1'b0;
                  active_thread[(149*4)+2] <= 1'b0;
                  active_thread[(149*4)+3] <= 1'b0;
                  spc149_inst_done         <= 0;
                  spc149_phy_pc_w          <= 0;
                end else begin
                  active_thread[(149*4)]   <= 1'b1;
                  active_thread[(149*4)+1] <= 1'b1;
                  active_thread[(149*4)+2] <= 1'b1;
                  active_thread[(149*4)+3] <= 1'b1;
                  spc149_inst_done         <= `ARIANE_CORE149.piton_pc_vld;
                  spc149_phy_pc_w          <= `ARIANE_CORE149.piton_pc;
                end
            end
    

            assign spc150_thread_id = 2'b00;
            assign spc150_rtl_pc = spc150_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(150*4)]   <= 1'b0;
                  active_thread[(150*4)+1] <= 1'b0;
                  active_thread[(150*4)+2] <= 1'b0;
                  active_thread[(150*4)+3] <= 1'b0;
                  spc150_inst_done         <= 0;
                  spc150_phy_pc_w          <= 0;
                end else begin
                  active_thread[(150*4)]   <= 1'b1;
                  active_thread[(150*4)+1] <= 1'b1;
                  active_thread[(150*4)+2] <= 1'b1;
                  active_thread[(150*4)+3] <= 1'b1;
                  spc150_inst_done         <= `ARIANE_CORE150.piton_pc_vld;
                  spc150_phy_pc_w          <= `ARIANE_CORE150.piton_pc;
                end
            end
    

            assign spc151_thread_id = 2'b00;
            assign spc151_rtl_pc = spc151_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(151*4)]   <= 1'b0;
                  active_thread[(151*4)+1] <= 1'b0;
                  active_thread[(151*4)+2] <= 1'b0;
                  active_thread[(151*4)+3] <= 1'b0;
                  spc151_inst_done         <= 0;
                  spc151_phy_pc_w          <= 0;
                end else begin
                  active_thread[(151*4)]   <= 1'b1;
                  active_thread[(151*4)+1] <= 1'b1;
                  active_thread[(151*4)+2] <= 1'b1;
                  active_thread[(151*4)+3] <= 1'b1;
                  spc151_inst_done         <= `ARIANE_CORE151.piton_pc_vld;
                  spc151_phy_pc_w          <= `ARIANE_CORE151.piton_pc;
                end
            end
    

            assign spc152_thread_id = 2'b00;
            assign spc152_rtl_pc = spc152_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(152*4)]   <= 1'b0;
                  active_thread[(152*4)+1] <= 1'b0;
                  active_thread[(152*4)+2] <= 1'b0;
                  active_thread[(152*4)+3] <= 1'b0;
                  spc152_inst_done         <= 0;
                  spc152_phy_pc_w          <= 0;
                end else begin
                  active_thread[(152*4)]   <= 1'b1;
                  active_thread[(152*4)+1] <= 1'b1;
                  active_thread[(152*4)+2] <= 1'b1;
                  active_thread[(152*4)+3] <= 1'b1;
                  spc152_inst_done         <= `ARIANE_CORE152.piton_pc_vld;
                  spc152_phy_pc_w          <= `ARIANE_CORE152.piton_pc;
                end
            end
    

            assign spc153_thread_id = 2'b00;
            assign spc153_rtl_pc = spc153_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(153*4)]   <= 1'b0;
                  active_thread[(153*4)+1] <= 1'b0;
                  active_thread[(153*4)+2] <= 1'b0;
                  active_thread[(153*4)+3] <= 1'b0;
                  spc153_inst_done         <= 0;
                  spc153_phy_pc_w          <= 0;
                end else begin
                  active_thread[(153*4)]   <= 1'b1;
                  active_thread[(153*4)+1] <= 1'b1;
                  active_thread[(153*4)+2] <= 1'b1;
                  active_thread[(153*4)+3] <= 1'b1;
                  spc153_inst_done         <= `ARIANE_CORE153.piton_pc_vld;
                  spc153_phy_pc_w          <= `ARIANE_CORE153.piton_pc;
                end
            end
    

            assign spc154_thread_id = 2'b00;
            assign spc154_rtl_pc = spc154_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(154*4)]   <= 1'b0;
                  active_thread[(154*4)+1] <= 1'b0;
                  active_thread[(154*4)+2] <= 1'b0;
                  active_thread[(154*4)+3] <= 1'b0;
                  spc154_inst_done         <= 0;
                  spc154_phy_pc_w          <= 0;
                end else begin
                  active_thread[(154*4)]   <= 1'b1;
                  active_thread[(154*4)+1] <= 1'b1;
                  active_thread[(154*4)+2] <= 1'b1;
                  active_thread[(154*4)+3] <= 1'b1;
                  spc154_inst_done         <= `ARIANE_CORE154.piton_pc_vld;
                  spc154_phy_pc_w          <= `ARIANE_CORE154.piton_pc;
                end
            end
    

            assign spc155_thread_id = 2'b00;
            assign spc155_rtl_pc = spc155_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(155*4)]   <= 1'b0;
                  active_thread[(155*4)+1] <= 1'b0;
                  active_thread[(155*4)+2] <= 1'b0;
                  active_thread[(155*4)+3] <= 1'b0;
                  spc155_inst_done         <= 0;
                  spc155_phy_pc_w          <= 0;
                end else begin
                  active_thread[(155*4)]   <= 1'b1;
                  active_thread[(155*4)+1] <= 1'b1;
                  active_thread[(155*4)+2] <= 1'b1;
                  active_thread[(155*4)+3] <= 1'b1;
                  spc155_inst_done         <= `ARIANE_CORE155.piton_pc_vld;
                  spc155_phy_pc_w          <= `ARIANE_CORE155.piton_pc;
                end
            end
    

            assign spc156_thread_id = 2'b00;
            assign spc156_rtl_pc = spc156_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(156*4)]   <= 1'b0;
                  active_thread[(156*4)+1] <= 1'b0;
                  active_thread[(156*4)+2] <= 1'b0;
                  active_thread[(156*4)+3] <= 1'b0;
                  spc156_inst_done         <= 0;
                  spc156_phy_pc_w          <= 0;
                end else begin
                  active_thread[(156*4)]   <= 1'b1;
                  active_thread[(156*4)+1] <= 1'b1;
                  active_thread[(156*4)+2] <= 1'b1;
                  active_thread[(156*4)+3] <= 1'b1;
                  spc156_inst_done         <= `ARIANE_CORE156.piton_pc_vld;
                  spc156_phy_pc_w          <= `ARIANE_CORE156.piton_pc;
                end
            end
    

            assign spc157_thread_id = 2'b00;
            assign spc157_rtl_pc = spc157_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(157*4)]   <= 1'b0;
                  active_thread[(157*4)+1] <= 1'b0;
                  active_thread[(157*4)+2] <= 1'b0;
                  active_thread[(157*4)+3] <= 1'b0;
                  spc157_inst_done         <= 0;
                  spc157_phy_pc_w          <= 0;
                end else begin
                  active_thread[(157*4)]   <= 1'b1;
                  active_thread[(157*4)+1] <= 1'b1;
                  active_thread[(157*4)+2] <= 1'b1;
                  active_thread[(157*4)+3] <= 1'b1;
                  spc157_inst_done         <= `ARIANE_CORE157.piton_pc_vld;
                  spc157_phy_pc_w          <= `ARIANE_CORE157.piton_pc;
                end
            end
    

            assign spc158_thread_id = 2'b00;
            assign spc158_rtl_pc = spc158_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(158*4)]   <= 1'b0;
                  active_thread[(158*4)+1] <= 1'b0;
                  active_thread[(158*4)+2] <= 1'b0;
                  active_thread[(158*4)+3] <= 1'b0;
                  spc158_inst_done         <= 0;
                  spc158_phy_pc_w          <= 0;
                end else begin
                  active_thread[(158*4)]   <= 1'b1;
                  active_thread[(158*4)+1] <= 1'b1;
                  active_thread[(158*4)+2] <= 1'b1;
                  active_thread[(158*4)+3] <= 1'b1;
                  spc158_inst_done         <= `ARIANE_CORE158.piton_pc_vld;
                  spc158_phy_pc_w          <= `ARIANE_CORE158.piton_pc;
                end
            end
    

            assign spc159_thread_id = 2'b00;
            assign spc159_rtl_pc = spc159_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(159*4)]   <= 1'b0;
                  active_thread[(159*4)+1] <= 1'b0;
                  active_thread[(159*4)+2] <= 1'b0;
                  active_thread[(159*4)+3] <= 1'b0;
                  spc159_inst_done         <= 0;
                  spc159_phy_pc_w          <= 0;
                end else begin
                  active_thread[(159*4)]   <= 1'b1;
                  active_thread[(159*4)+1] <= 1'b1;
                  active_thread[(159*4)+2] <= 1'b1;
                  active_thread[(159*4)+3] <= 1'b1;
                  spc159_inst_done         <= `ARIANE_CORE159.piton_pc_vld;
                  spc159_phy_pc_w          <= `ARIANE_CORE159.piton_pc;
                end
            end
    

            assign spc160_thread_id = 2'b00;
            assign spc160_rtl_pc = spc160_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(160*4)]   <= 1'b0;
                  active_thread[(160*4)+1] <= 1'b0;
                  active_thread[(160*4)+2] <= 1'b0;
                  active_thread[(160*4)+3] <= 1'b0;
                  spc160_inst_done         <= 0;
                  spc160_phy_pc_w          <= 0;
                end else begin
                  active_thread[(160*4)]   <= 1'b1;
                  active_thread[(160*4)+1] <= 1'b1;
                  active_thread[(160*4)+2] <= 1'b1;
                  active_thread[(160*4)+3] <= 1'b1;
                  spc160_inst_done         <= `ARIANE_CORE160.piton_pc_vld;
                  spc160_phy_pc_w          <= `ARIANE_CORE160.piton_pc;
                end
            end
    

            assign spc161_thread_id = 2'b00;
            assign spc161_rtl_pc = spc161_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(161*4)]   <= 1'b0;
                  active_thread[(161*4)+1] <= 1'b0;
                  active_thread[(161*4)+2] <= 1'b0;
                  active_thread[(161*4)+3] <= 1'b0;
                  spc161_inst_done         <= 0;
                  spc161_phy_pc_w          <= 0;
                end else begin
                  active_thread[(161*4)]   <= 1'b1;
                  active_thread[(161*4)+1] <= 1'b1;
                  active_thread[(161*4)+2] <= 1'b1;
                  active_thread[(161*4)+3] <= 1'b1;
                  spc161_inst_done         <= `ARIANE_CORE161.piton_pc_vld;
                  spc161_phy_pc_w          <= `ARIANE_CORE161.piton_pc;
                end
            end
    

            assign spc162_thread_id = 2'b00;
            assign spc162_rtl_pc = spc162_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(162*4)]   <= 1'b0;
                  active_thread[(162*4)+1] <= 1'b0;
                  active_thread[(162*4)+2] <= 1'b0;
                  active_thread[(162*4)+3] <= 1'b0;
                  spc162_inst_done         <= 0;
                  spc162_phy_pc_w          <= 0;
                end else begin
                  active_thread[(162*4)]   <= 1'b1;
                  active_thread[(162*4)+1] <= 1'b1;
                  active_thread[(162*4)+2] <= 1'b1;
                  active_thread[(162*4)+3] <= 1'b1;
                  spc162_inst_done         <= `ARIANE_CORE162.piton_pc_vld;
                  spc162_phy_pc_w          <= `ARIANE_CORE162.piton_pc;
                end
            end
    

            assign spc163_thread_id = 2'b00;
            assign spc163_rtl_pc = spc163_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(163*4)]   <= 1'b0;
                  active_thread[(163*4)+1] <= 1'b0;
                  active_thread[(163*4)+2] <= 1'b0;
                  active_thread[(163*4)+3] <= 1'b0;
                  spc163_inst_done         <= 0;
                  spc163_phy_pc_w          <= 0;
                end else begin
                  active_thread[(163*4)]   <= 1'b1;
                  active_thread[(163*4)+1] <= 1'b1;
                  active_thread[(163*4)+2] <= 1'b1;
                  active_thread[(163*4)+3] <= 1'b1;
                  spc163_inst_done         <= `ARIANE_CORE163.piton_pc_vld;
                  spc163_phy_pc_w          <= `ARIANE_CORE163.piton_pc;
                end
            end
    

            assign spc164_thread_id = 2'b00;
            assign spc164_rtl_pc = spc164_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(164*4)]   <= 1'b0;
                  active_thread[(164*4)+1] <= 1'b0;
                  active_thread[(164*4)+2] <= 1'b0;
                  active_thread[(164*4)+3] <= 1'b0;
                  spc164_inst_done         <= 0;
                  spc164_phy_pc_w          <= 0;
                end else begin
                  active_thread[(164*4)]   <= 1'b1;
                  active_thread[(164*4)+1] <= 1'b1;
                  active_thread[(164*4)+2] <= 1'b1;
                  active_thread[(164*4)+3] <= 1'b1;
                  spc164_inst_done         <= `ARIANE_CORE164.piton_pc_vld;
                  spc164_phy_pc_w          <= `ARIANE_CORE164.piton_pc;
                end
            end
    

            assign spc165_thread_id = 2'b00;
            assign spc165_rtl_pc = spc165_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(165*4)]   <= 1'b0;
                  active_thread[(165*4)+1] <= 1'b0;
                  active_thread[(165*4)+2] <= 1'b0;
                  active_thread[(165*4)+3] <= 1'b0;
                  spc165_inst_done         <= 0;
                  spc165_phy_pc_w          <= 0;
                end else begin
                  active_thread[(165*4)]   <= 1'b1;
                  active_thread[(165*4)+1] <= 1'b1;
                  active_thread[(165*4)+2] <= 1'b1;
                  active_thread[(165*4)+3] <= 1'b1;
                  spc165_inst_done         <= `ARIANE_CORE165.piton_pc_vld;
                  spc165_phy_pc_w          <= `ARIANE_CORE165.piton_pc;
                end
            end
    

            assign spc166_thread_id = 2'b00;
            assign spc166_rtl_pc = spc166_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(166*4)]   <= 1'b0;
                  active_thread[(166*4)+1] <= 1'b0;
                  active_thread[(166*4)+2] <= 1'b0;
                  active_thread[(166*4)+3] <= 1'b0;
                  spc166_inst_done         <= 0;
                  spc166_phy_pc_w          <= 0;
                end else begin
                  active_thread[(166*4)]   <= 1'b1;
                  active_thread[(166*4)+1] <= 1'b1;
                  active_thread[(166*4)+2] <= 1'b1;
                  active_thread[(166*4)+3] <= 1'b1;
                  spc166_inst_done         <= `ARIANE_CORE166.piton_pc_vld;
                  spc166_phy_pc_w          <= `ARIANE_CORE166.piton_pc;
                end
            end
    

            assign spc167_thread_id = 2'b00;
            assign spc167_rtl_pc = spc167_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(167*4)]   <= 1'b0;
                  active_thread[(167*4)+1] <= 1'b0;
                  active_thread[(167*4)+2] <= 1'b0;
                  active_thread[(167*4)+3] <= 1'b0;
                  spc167_inst_done         <= 0;
                  spc167_phy_pc_w          <= 0;
                end else begin
                  active_thread[(167*4)]   <= 1'b1;
                  active_thread[(167*4)+1] <= 1'b1;
                  active_thread[(167*4)+2] <= 1'b1;
                  active_thread[(167*4)+3] <= 1'b1;
                  spc167_inst_done         <= `ARIANE_CORE167.piton_pc_vld;
                  spc167_phy_pc_w          <= `ARIANE_CORE167.piton_pc;
                end
            end
    

            assign spc168_thread_id = 2'b00;
            assign spc168_rtl_pc = spc168_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(168*4)]   <= 1'b0;
                  active_thread[(168*4)+1] <= 1'b0;
                  active_thread[(168*4)+2] <= 1'b0;
                  active_thread[(168*4)+3] <= 1'b0;
                  spc168_inst_done         <= 0;
                  spc168_phy_pc_w          <= 0;
                end else begin
                  active_thread[(168*4)]   <= 1'b1;
                  active_thread[(168*4)+1] <= 1'b1;
                  active_thread[(168*4)+2] <= 1'b1;
                  active_thread[(168*4)+3] <= 1'b1;
                  spc168_inst_done         <= `ARIANE_CORE168.piton_pc_vld;
                  spc168_phy_pc_w          <= `ARIANE_CORE168.piton_pc;
                end
            end
    

            assign spc169_thread_id = 2'b00;
            assign spc169_rtl_pc = spc169_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(169*4)]   <= 1'b0;
                  active_thread[(169*4)+1] <= 1'b0;
                  active_thread[(169*4)+2] <= 1'b0;
                  active_thread[(169*4)+3] <= 1'b0;
                  spc169_inst_done         <= 0;
                  spc169_phy_pc_w          <= 0;
                end else begin
                  active_thread[(169*4)]   <= 1'b1;
                  active_thread[(169*4)+1] <= 1'b1;
                  active_thread[(169*4)+2] <= 1'b1;
                  active_thread[(169*4)+3] <= 1'b1;
                  spc169_inst_done         <= `ARIANE_CORE169.piton_pc_vld;
                  spc169_phy_pc_w          <= `ARIANE_CORE169.piton_pc;
                end
            end
    

            assign spc170_thread_id = 2'b00;
            assign spc170_rtl_pc = spc170_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(170*4)]   <= 1'b0;
                  active_thread[(170*4)+1] <= 1'b0;
                  active_thread[(170*4)+2] <= 1'b0;
                  active_thread[(170*4)+3] <= 1'b0;
                  spc170_inst_done         <= 0;
                  spc170_phy_pc_w          <= 0;
                end else begin
                  active_thread[(170*4)]   <= 1'b1;
                  active_thread[(170*4)+1] <= 1'b1;
                  active_thread[(170*4)+2] <= 1'b1;
                  active_thread[(170*4)+3] <= 1'b1;
                  spc170_inst_done         <= `ARIANE_CORE170.piton_pc_vld;
                  spc170_phy_pc_w          <= `ARIANE_CORE170.piton_pc;
                end
            end
    

            assign spc171_thread_id = 2'b00;
            assign spc171_rtl_pc = spc171_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(171*4)]   <= 1'b0;
                  active_thread[(171*4)+1] <= 1'b0;
                  active_thread[(171*4)+2] <= 1'b0;
                  active_thread[(171*4)+3] <= 1'b0;
                  spc171_inst_done         <= 0;
                  spc171_phy_pc_w          <= 0;
                end else begin
                  active_thread[(171*4)]   <= 1'b1;
                  active_thread[(171*4)+1] <= 1'b1;
                  active_thread[(171*4)+2] <= 1'b1;
                  active_thread[(171*4)+3] <= 1'b1;
                  spc171_inst_done         <= `ARIANE_CORE171.piton_pc_vld;
                  spc171_phy_pc_w          <= `ARIANE_CORE171.piton_pc;
                end
            end
    

            assign spc172_thread_id = 2'b00;
            assign spc172_rtl_pc = spc172_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(172*4)]   <= 1'b0;
                  active_thread[(172*4)+1] <= 1'b0;
                  active_thread[(172*4)+2] <= 1'b0;
                  active_thread[(172*4)+3] <= 1'b0;
                  spc172_inst_done         <= 0;
                  spc172_phy_pc_w          <= 0;
                end else begin
                  active_thread[(172*4)]   <= 1'b1;
                  active_thread[(172*4)+1] <= 1'b1;
                  active_thread[(172*4)+2] <= 1'b1;
                  active_thread[(172*4)+3] <= 1'b1;
                  spc172_inst_done         <= `ARIANE_CORE172.piton_pc_vld;
                  spc172_phy_pc_w          <= `ARIANE_CORE172.piton_pc;
                end
            end
    

            assign spc173_thread_id = 2'b00;
            assign spc173_rtl_pc = spc173_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(173*4)]   <= 1'b0;
                  active_thread[(173*4)+1] <= 1'b0;
                  active_thread[(173*4)+2] <= 1'b0;
                  active_thread[(173*4)+3] <= 1'b0;
                  spc173_inst_done         <= 0;
                  spc173_phy_pc_w          <= 0;
                end else begin
                  active_thread[(173*4)]   <= 1'b1;
                  active_thread[(173*4)+1] <= 1'b1;
                  active_thread[(173*4)+2] <= 1'b1;
                  active_thread[(173*4)+3] <= 1'b1;
                  spc173_inst_done         <= `ARIANE_CORE173.piton_pc_vld;
                  spc173_phy_pc_w          <= `ARIANE_CORE173.piton_pc;
                end
            end
    

            assign spc174_thread_id = 2'b00;
            assign spc174_rtl_pc = spc174_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(174*4)]   <= 1'b0;
                  active_thread[(174*4)+1] <= 1'b0;
                  active_thread[(174*4)+2] <= 1'b0;
                  active_thread[(174*4)+3] <= 1'b0;
                  spc174_inst_done         <= 0;
                  spc174_phy_pc_w          <= 0;
                end else begin
                  active_thread[(174*4)]   <= 1'b1;
                  active_thread[(174*4)+1] <= 1'b1;
                  active_thread[(174*4)+2] <= 1'b1;
                  active_thread[(174*4)+3] <= 1'b1;
                  spc174_inst_done         <= `ARIANE_CORE174.piton_pc_vld;
                  spc174_phy_pc_w          <= `ARIANE_CORE174.piton_pc;
                end
            end
    

            assign spc175_thread_id = 2'b00;
            assign spc175_rtl_pc = spc175_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(175*4)]   <= 1'b0;
                  active_thread[(175*4)+1] <= 1'b0;
                  active_thread[(175*4)+2] <= 1'b0;
                  active_thread[(175*4)+3] <= 1'b0;
                  spc175_inst_done         <= 0;
                  spc175_phy_pc_w          <= 0;
                end else begin
                  active_thread[(175*4)]   <= 1'b1;
                  active_thread[(175*4)+1] <= 1'b1;
                  active_thread[(175*4)+2] <= 1'b1;
                  active_thread[(175*4)+3] <= 1'b1;
                  spc175_inst_done         <= `ARIANE_CORE175.piton_pc_vld;
                  spc175_phy_pc_w          <= `ARIANE_CORE175.piton_pc;
                end
            end
    

            assign spc176_thread_id = 2'b00;
            assign spc176_rtl_pc = spc176_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(176*4)]   <= 1'b0;
                  active_thread[(176*4)+1] <= 1'b0;
                  active_thread[(176*4)+2] <= 1'b0;
                  active_thread[(176*4)+3] <= 1'b0;
                  spc176_inst_done         <= 0;
                  spc176_phy_pc_w          <= 0;
                end else begin
                  active_thread[(176*4)]   <= 1'b1;
                  active_thread[(176*4)+1] <= 1'b1;
                  active_thread[(176*4)+2] <= 1'b1;
                  active_thread[(176*4)+3] <= 1'b1;
                  spc176_inst_done         <= `ARIANE_CORE176.piton_pc_vld;
                  spc176_phy_pc_w          <= `ARIANE_CORE176.piton_pc;
                end
            end
    

            assign spc177_thread_id = 2'b00;
            assign spc177_rtl_pc = spc177_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(177*4)]   <= 1'b0;
                  active_thread[(177*4)+1] <= 1'b0;
                  active_thread[(177*4)+2] <= 1'b0;
                  active_thread[(177*4)+3] <= 1'b0;
                  spc177_inst_done         <= 0;
                  spc177_phy_pc_w          <= 0;
                end else begin
                  active_thread[(177*4)]   <= 1'b1;
                  active_thread[(177*4)+1] <= 1'b1;
                  active_thread[(177*4)+2] <= 1'b1;
                  active_thread[(177*4)+3] <= 1'b1;
                  spc177_inst_done         <= `ARIANE_CORE177.piton_pc_vld;
                  spc177_phy_pc_w          <= `ARIANE_CORE177.piton_pc;
                end
            end
    

            assign spc178_thread_id = 2'b00;
            assign spc178_rtl_pc = spc178_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(178*4)]   <= 1'b0;
                  active_thread[(178*4)+1] <= 1'b0;
                  active_thread[(178*4)+2] <= 1'b0;
                  active_thread[(178*4)+3] <= 1'b0;
                  spc178_inst_done         <= 0;
                  spc178_phy_pc_w          <= 0;
                end else begin
                  active_thread[(178*4)]   <= 1'b1;
                  active_thread[(178*4)+1] <= 1'b1;
                  active_thread[(178*4)+2] <= 1'b1;
                  active_thread[(178*4)+3] <= 1'b1;
                  spc178_inst_done         <= `ARIANE_CORE178.piton_pc_vld;
                  spc178_phy_pc_w          <= `ARIANE_CORE178.piton_pc;
                end
            end
    

            assign spc179_thread_id = 2'b00;
            assign spc179_rtl_pc = spc179_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(179*4)]   <= 1'b0;
                  active_thread[(179*4)+1] <= 1'b0;
                  active_thread[(179*4)+2] <= 1'b0;
                  active_thread[(179*4)+3] <= 1'b0;
                  spc179_inst_done         <= 0;
                  spc179_phy_pc_w          <= 0;
                end else begin
                  active_thread[(179*4)]   <= 1'b1;
                  active_thread[(179*4)+1] <= 1'b1;
                  active_thread[(179*4)+2] <= 1'b1;
                  active_thread[(179*4)+3] <= 1'b1;
                  spc179_inst_done         <= `ARIANE_CORE179.piton_pc_vld;
                  spc179_phy_pc_w          <= `ARIANE_CORE179.piton_pc;
                end
            end
    

            assign spc180_thread_id = 2'b00;
            assign spc180_rtl_pc = spc180_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(180*4)]   <= 1'b0;
                  active_thread[(180*4)+1] <= 1'b0;
                  active_thread[(180*4)+2] <= 1'b0;
                  active_thread[(180*4)+3] <= 1'b0;
                  spc180_inst_done         <= 0;
                  spc180_phy_pc_w          <= 0;
                end else begin
                  active_thread[(180*4)]   <= 1'b1;
                  active_thread[(180*4)+1] <= 1'b1;
                  active_thread[(180*4)+2] <= 1'b1;
                  active_thread[(180*4)+3] <= 1'b1;
                  spc180_inst_done         <= `ARIANE_CORE180.piton_pc_vld;
                  spc180_phy_pc_w          <= `ARIANE_CORE180.piton_pc;
                end
            end
    

            assign spc181_thread_id = 2'b00;
            assign spc181_rtl_pc = spc181_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(181*4)]   <= 1'b0;
                  active_thread[(181*4)+1] <= 1'b0;
                  active_thread[(181*4)+2] <= 1'b0;
                  active_thread[(181*4)+3] <= 1'b0;
                  spc181_inst_done         <= 0;
                  spc181_phy_pc_w          <= 0;
                end else begin
                  active_thread[(181*4)]   <= 1'b1;
                  active_thread[(181*4)+1] <= 1'b1;
                  active_thread[(181*4)+2] <= 1'b1;
                  active_thread[(181*4)+3] <= 1'b1;
                  spc181_inst_done         <= `ARIANE_CORE181.piton_pc_vld;
                  spc181_phy_pc_w          <= `ARIANE_CORE181.piton_pc;
                end
            end
    

            assign spc182_thread_id = 2'b00;
            assign spc182_rtl_pc = spc182_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(182*4)]   <= 1'b0;
                  active_thread[(182*4)+1] <= 1'b0;
                  active_thread[(182*4)+2] <= 1'b0;
                  active_thread[(182*4)+3] <= 1'b0;
                  spc182_inst_done         <= 0;
                  spc182_phy_pc_w          <= 0;
                end else begin
                  active_thread[(182*4)]   <= 1'b1;
                  active_thread[(182*4)+1] <= 1'b1;
                  active_thread[(182*4)+2] <= 1'b1;
                  active_thread[(182*4)+3] <= 1'b1;
                  spc182_inst_done         <= `ARIANE_CORE182.piton_pc_vld;
                  spc182_phy_pc_w          <= `ARIANE_CORE182.piton_pc;
                end
            end
    

            assign spc183_thread_id = 2'b00;
            assign spc183_rtl_pc = spc183_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(183*4)]   <= 1'b0;
                  active_thread[(183*4)+1] <= 1'b0;
                  active_thread[(183*4)+2] <= 1'b0;
                  active_thread[(183*4)+3] <= 1'b0;
                  spc183_inst_done         <= 0;
                  spc183_phy_pc_w          <= 0;
                end else begin
                  active_thread[(183*4)]   <= 1'b1;
                  active_thread[(183*4)+1] <= 1'b1;
                  active_thread[(183*4)+2] <= 1'b1;
                  active_thread[(183*4)+3] <= 1'b1;
                  spc183_inst_done         <= `ARIANE_CORE183.piton_pc_vld;
                  spc183_phy_pc_w          <= `ARIANE_CORE183.piton_pc;
                end
            end
    

            assign spc184_thread_id = 2'b00;
            assign spc184_rtl_pc = spc184_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(184*4)]   <= 1'b0;
                  active_thread[(184*4)+1] <= 1'b0;
                  active_thread[(184*4)+2] <= 1'b0;
                  active_thread[(184*4)+3] <= 1'b0;
                  spc184_inst_done         <= 0;
                  spc184_phy_pc_w          <= 0;
                end else begin
                  active_thread[(184*4)]   <= 1'b1;
                  active_thread[(184*4)+1] <= 1'b1;
                  active_thread[(184*4)+2] <= 1'b1;
                  active_thread[(184*4)+3] <= 1'b1;
                  spc184_inst_done         <= `ARIANE_CORE184.piton_pc_vld;
                  spc184_phy_pc_w          <= `ARIANE_CORE184.piton_pc;
                end
            end
    

            assign spc185_thread_id = 2'b00;
            assign spc185_rtl_pc = spc185_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(185*4)]   <= 1'b0;
                  active_thread[(185*4)+1] <= 1'b0;
                  active_thread[(185*4)+2] <= 1'b0;
                  active_thread[(185*4)+3] <= 1'b0;
                  spc185_inst_done         <= 0;
                  spc185_phy_pc_w          <= 0;
                end else begin
                  active_thread[(185*4)]   <= 1'b1;
                  active_thread[(185*4)+1] <= 1'b1;
                  active_thread[(185*4)+2] <= 1'b1;
                  active_thread[(185*4)+3] <= 1'b1;
                  spc185_inst_done         <= `ARIANE_CORE185.piton_pc_vld;
                  spc185_phy_pc_w          <= `ARIANE_CORE185.piton_pc;
                end
            end
    

            assign spc186_thread_id = 2'b00;
            assign spc186_rtl_pc = spc186_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(186*4)]   <= 1'b0;
                  active_thread[(186*4)+1] <= 1'b0;
                  active_thread[(186*4)+2] <= 1'b0;
                  active_thread[(186*4)+3] <= 1'b0;
                  spc186_inst_done         <= 0;
                  spc186_phy_pc_w          <= 0;
                end else begin
                  active_thread[(186*4)]   <= 1'b1;
                  active_thread[(186*4)+1] <= 1'b1;
                  active_thread[(186*4)+2] <= 1'b1;
                  active_thread[(186*4)+3] <= 1'b1;
                  spc186_inst_done         <= `ARIANE_CORE186.piton_pc_vld;
                  spc186_phy_pc_w          <= `ARIANE_CORE186.piton_pc;
                end
            end
    

            assign spc187_thread_id = 2'b00;
            assign spc187_rtl_pc = spc187_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(187*4)]   <= 1'b0;
                  active_thread[(187*4)+1] <= 1'b0;
                  active_thread[(187*4)+2] <= 1'b0;
                  active_thread[(187*4)+3] <= 1'b0;
                  spc187_inst_done         <= 0;
                  spc187_phy_pc_w          <= 0;
                end else begin
                  active_thread[(187*4)]   <= 1'b1;
                  active_thread[(187*4)+1] <= 1'b1;
                  active_thread[(187*4)+2] <= 1'b1;
                  active_thread[(187*4)+3] <= 1'b1;
                  spc187_inst_done         <= `ARIANE_CORE187.piton_pc_vld;
                  spc187_phy_pc_w          <= `ARIANE_CORE187.piton_pc;
                end
            end
    

            assign spc188_thread_id = 2'b00;
            assign spc188_rtl_pc = spc188_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(188*4)]   <= 1'b0;
                  active_thread[(188*4)+1] <= 1'b0;
                  active_thread[(188*4)+2] <= 1'b0;
                  active_thread[(188*4)+3] <= 1'b0;
                  spc188_inst_done         <= 0;
                  spc188_phy_pc_w          <= 0;
                end else begin
                  active_thread[(188*4)]   <= 1'b1;
                  active_thread[(188*4)+1] <= 1'b1;
                  active_thread[(188*4)+2] <= 1'b1;
                  active_thread[(188*4)+3] <= 1'b1;
                  spc188_inst_done         <= `ARIANE_CORE188.piton_pc_vld;
                  spc188_phy_pc_w          <= `ARIANE_CORE188.piton_pc;
                end
            end
    

            assign spc189_thread_id = 2'b00;
            assign spc189_rtl_pc = spc189_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(189*4)]   <= 1'b0;
                  active_thread[(189*4)+1] <= 1'b0;
                  active_thread[(189*4)+2] <= 1'b0;
                  active_thread[(189*4)+3] <= 1'b0;
                  spc189_inst_done         <= 0;
                  spc189_phy_pc_w          <= 0;
                end else begin
                  active_thread[(189*4)]   <= 1'b1;
                  active_thread[(189*4)+1] <= 1'b1;
                  active_thread[(189*4)+2] <= 1'b1;
                  active_thread[(189*4)+3] <= 1'b1;
                  spc189_inst_done         <= `ARIANE_CORE189.piton_pc_vld;
                  spc189_phy_pc_w          <= `ARIANE_CORE189.piton_pc;
                end
            end
    

            assign spc190_thread_id = 2'b00;
            assign spc190_rtl_pc = spc190_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(190*4)]   <= 1'b0;
                  active_thread[(190*4)+1] <= 1'b0;
                  active_thread[(190*4)+2] <= 1'b0;
                  active_thread[(190*4)+3] <= 1'b0;
                  spc190_inst_done         <= 0;
                  spc190_phy_pc_w          <= 0;
                end else begin
                  active_thread[(190*4)]   <= 1'b1;
                  active_thread[(190*4)+1] <= 1'b1;
                  active_thread[(190*4)+2] <= 1'b1;
                  active_thread[(190*4)+3] <= 1'b1;
                  spc190_inst_done         <= `ARIANE_CORE190.piton_pc_vld;
                  spc190_phy_pc_w          <= `ARIANE_CORE190.piton_pc;
                end
            end
    

            assign spc191_thread_id = 2'b00;
            assign spc191_rtl_pc = spc191_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(191*4)]   <= 1'b0;
                  active_thread[(191*4)+1] <= 1'b0;
                  active_thread[(191*4)+2] <= 1'b0;
                  active_thread[(191*4)+3] <= 1'b0;
                  spc191_inst_done         <= 0;
                  spc191_phy_pc_w          <= 0;
                end else begin
                  active_thread[(191*4)]   <= 1'b1;
                  active_thread[(191*4)+1] <= 1'b1;
                  active_thread[(191*4)+2] <= 1'b1;
                  active_thread[(191*4)+3] <= 1'b1;
                  spc191_inst_done         <= `ARIANE_CORE191.piton_pc_vld;
                  spc191_phy_pc_w          <= `ARIANE_CORE191.piton_pc;
                end
            end
    

            assign spc192_thread_id = 2'b00;
            assign spc192_rtl_pc = spc192_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(192*4)]   <= 1'b0;
                  active_thread[(192*4)+1] <= 1'b0;
                  active_thread[(192*4)+2] <= 1'b0;
                  active_thread[(192*4)+3] <= 1'b0;
                  spc192_inst_done         <= 0;
                  spc192_phy_pc_w          <= 0;
                end else begin
                  active_thread[(192*4)]   <= 1'b1;
                  active_thread[(192*4)+1] <= 1'b1;
                  active_thread[(192*4)+2] <= 1'b1;
                  active_thread[(192*4)+3] <= 1'b1;
                  spc192_inst_done         <= `ARIANE_CORE192.piton_pc_vld;
                  spc192_phy_pc_w          <= `ARIANE_CORE192.piton_pc;
                end
            end
    

            assign spc193_thread_id = 2'b00;
            assign spc193_rtl_pc = spc193_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(193*4)]   <= 1'b0;
                  active_thread[(193*4)+1] <= 1'b0;
                  active_thread[(193*4)+2] <= 1'b0;
                  active_thread[(193*4)+3] <= 1'b0;
                  spc193_inst_done         <= 0;
                  spc193_phy_pc_w          <= 0;
                end else begin
                  active_thread[(193*4)]   <= 1'b1;
                  active_thread[(193*4)+1] <= 1'b1;
                  active_thread[(193*4)+2] <= 1'b1;
                  active_thread[(193*4)+3] <= 1'b1;
                  spc193_inst_done         <= `ARIANE_CORE193.piton_pc_vld;
                  spc193_phy_pc_w          <= `ARIANE_CORE193.piton_pc;
                end
            end
    

            assign spc194_thread_id = 2'b00;
            assign spc194_rtl_pc = spc194_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(194*4)]   <= 1'b0;
                  active_thread[(194*4)+1] <= 1'b0;
                  active_thread[(194*4)+2] <= 1'b0;
                  active_thread[(194*4)+3] <= 1'b0;
                  spc194_inst_done         <= 0;
                  spc194_phy_pc_w          <= 0;
                end else begin
                  active_thread[(194*4)]   <= 1'b1;
                  active_thread[(194*4)+1] <= 1'b1;
                  active_thread[(194*4)+2] <= 1'b1;
                  active_thread[(194*4)+3] <= 1'b1;
                  spc194_inst_done         <= `ARIANE_CORE194.piton_pc_vld;
                  spc194_phy_pc_w          <= `ARIANE_CORE194.piton_pc;
                end
            end
    

            assign spc195_thread_id = 2'b00;
            assign spc195_rtl_pc = spc195_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(195*4)]   <= 1'b0;
                  active_thread[(195*4)+1] <= 1'b0;
                  active_thread[(195*4)+2] <= 1'b0;
                  active_thread[(195*4)+3] <= 1'b0;
                  spc195_inst_done         <= 0;
                  spc195_phy_pc_w          <= 0;
                end else begin
                  active_thread[(195*4)]   <= 1'b1;
                  active_thread[(195*4)+1] <= 1'b1;
                  active_thread[(195*4)+2] <= 1'b1;
                  active_thread[(195*4)+3] <= 1'b1;
                  spc195_inst_done         <= `ARIANE_CORE195.piton_pc_vld;
                  spc195_phy_pc_w          <= `ARIANE_CORE195.piton_pc;
                end
            end
    

            assign spc196_thread_id = 2'b00;
            assign spc196_rtl_pc = spc196_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(196*4)]   <= 1'b0;
                  active_thread[(196*4)+1] <= 1'b0;
                  active_thread[(196*4)+2] <= 1'b0;
                  active_thread[(196*4)+3] <= 1'b0;
                  spc196_inst_done         <= 0;
                  spc196_phy_pc_w          <= 0;
                end else begin
                  active_thread[(196*4)]   <= 1'b1;
                  active_thread[(196*4)+1] <= 1'b1;
                  active_thread[(196*4)+2] <= 1'b1;
                  active_thread[(196*4)+3] <= 1'b1;
                  spc196_inst_done         <= `ARIANE_CORE196.piton_pc_vld;
                  spc196_phy_pc_w          <= `ARIANE_CORE196.piton_pc;
                end
            end
    

            assign spc197_thread_id = 2'b00;
            assign spc197_rtl_pc = spc197_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(197*4)]   <= 1'b0;
                  active_thread[(197*4)+1] <= 1'b0;
                  active_thread[(197*4)+2] <= 1'b0;
                  active_thread[(197*4)+3] <= 1'b0;
                  spc197_inst_done         <= 0;
                  spc197_phy_pc_w          <= 0;
                end else begin
                  active_thread[(197*4)]   <= 1'b1;
                  active_thread[(197*4)+1] <= 1'b1;
                  active_thread[(197*4)+2] <= 1'b1;
                  active_thread[(197*4)+3] <= 1'b1;
                  spc197_inst_done         <= `ARIANE_CORE197.piton_pc_vld;
                  spc197_phy_pc_w          <= `ARIANE_CORE197.piton_pc;
                end
            end
    

            assign spc198_thread_id = 2'b00;
            assign spc198_rtl_pc = spc198_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(198*4)]   <= 1'b0;
                  active_thread[(198*4)+1] <= 1'b0;
                  active_thread[(198*4)+2] <= 1'b0;
                  active_thread[(198*4)+3] <= 1'b0;
                  spc198_inst_done         <= 0;
                  spc198_phy_pc_w          <= 0;
                end else begin
                  active_thread[(198*4)]   <= 1'b1;
                  active_thread[(198*4)+1] <= 1'b1;
                  active_thread[(198*4)+2] <= 1'b1;
                  active_thread[(198*4)+3] <= 1'b1;
                  spc198_inst_done         <= `ARIANE_CORE198.piton_pc_vld;
                  spc198_phy_pc_w          <= `ARIANE_CORE198.piton_pc;
                end
            end
    

            assign spc199_thread_id = 2'b00;
            assign spc199_rtl_pc = spc199_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(199*4)]   <= 1'b0;
                  active_thread[(199*4)+1] <= 1'b0;
                  active_thread[(199*4)+2] <= 1'b0;
                  active_thread[(199*4)+3] <= 1'b0;
                  spc199_inst_done         <= 0;
                  spc199_phy_pc_w          <= 0;
                end else begin
                  active_thread[(199*4)]   <= 1'b1;
                  active_thread[(199*4)+1] <= 1'b1;
                  active_thread[(199*4)+2] <= 1'b1;
                  active_thread[(199*4)+3] <= 1'b1;
                  spc199_inst_done         <= `ARIANE_CORE199.piton_pc_vld;
                  spc199_phy_pc_w          <= `ARIANE_CORE199.piton_pc;
                end
            end
    

            assign spc200_thread_id = 2'b00;
            assign spc200_rtl_pc = spc200_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(200*4)]   <= 1'b0;
                  active_thread[(200*4)+1] <= 1'b0;
                  active_thread[(200*4)+2] <= 1'b0;
                  active_thread[(200*4)+3] <= 1'b0;
                  spc200_inst_done         <= 0;
                  spc200_phy_pc_w          <= 0;
                end else begin
                  active_thread[(200*4)]   <= 1'b1;
                  active_thread[(200*4)+1] <= 1'b1;
                  active_thread[(200*4)+2] <= 1'b1;
                  active_thread[(200*4)+3] <= 1'b1;
                  spc200_inst_done         <= `ARIANE_CORE200.piton_pc_vld;
                  spc200_phy_pc_w          <= `ARIANE_CORE200.piton_pc;
                end
            end
    

            assign spc201_thread_id = 2'b00;
            assign spc201_rtl_pc = spc201_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(201*4)]   <= 1'b0;
                  active_thread[(201*4)+1] <= 1'b0;
                  active_thread[(201*4)+2] <= 1'b0;
                  active_thread[(201*4)+3] <= 1'b0;
                  spc201_inst_done         <= 0;
                  spc201_phy_pc_w          <= 0;
                end else begin
                  active_thread[(201*4)]   <= 1'b1;
                  active_thread[(201*4)+1] <= 1'b1;
                  active_thread[(201*4)+2] <= 1'b1;
                  active_thread[(201*4)+3] <= 1'b1;
                  spc201_inst_done         <= `ARIANE_CORE201.piton_pc_vld;
                  spc201_phy_pc_w          <= `ARIANE_CORE201.piton_pc;
                end
            end
    

            assign spc202_thread_id = 2'b00;
            assign spc202_rtl_pc = spc202_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(202*4)]   <= 1'b0;
                  active_thread[(202*4)+1] <= 1'b0;
                  active_thread[(202*4)+2] <= 1'b0;
                  active_thread[(202*4)+3] <= 1'b0;
                  spc202_inst_done         <= 0;
                  spc202_phy_pc_w          <= 0;
                end else begin
                  active_thread[(202*4)]   <= 1'b1;
                  active_thread[(202*4)+1] <= 1'b1;
                  active_thread[(202*4)+2] <= 1'b1;
                  active_thread[(202*4)+3] <= 1'b1;
                  spc202_inst_done         <= `ARIANE_CORE202.piton_pc_vld;
                  spc202_phy_pc_w          <= `ARIANE_CORE202.piton_pc;
                end
            end
    

            assign spc203_thread_id = 2'b00;
            assign spc203_rtl_pc = spc203_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(203*4)]   <= 1'b0;
                  active_thread[(203*4)+1] <= 1'b0;
                  active_thread[(203*4)+2] <= 1'b0;
                  active_thread[(203*4)+3] <= 1'b0;
                  spc203_inst_done         <= 0;
                  spc203_phy_pc_w          <= 0;
                end else begin
                  active_thread[(203*4)]   <= 1'b1;
                  active_thread[(203*4)+1] <= 1'b1;
                  active_thread[(203*4)+2] <= 1'b1;
                  active_thread[(203*4)+3] <= 1'b1;
                  spc203_inst_done         <= `ARIANE_CORE203.piton_pc_vld;
                  spc203_phy_pc_w          <= `ARIANE_CORE203.piton_pc;
                end
            end
    

            assign spc204_thread_id = 2'b00;
            assign spc204_rtl_pc = spc204_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(204*4)]   <= 1'b0;
                  active_thread[(204*4)+1] <= 1'b0;
                  active_thread[(204*4)+2] <= 1'b0;
                  active_thread[(204*4)+3] <= 1'b0;
                  spc204_inst_done         <= 0;
                  spc204_phy_pc_w          <= 0;
                end else begin
                  active_thread[(204*4)]   <= 1'b1;
                  active_thread[(204*4)+1] <= 1'b1;
                  active_thread[(204*4)+2] <= 1'b1;
                  active_thread[(204*4)+3] <= 1'b1;
                  spc204_inst_done         <= `ARIANE_CORE204.piton_pc_vld;
                  spc204_phy_pc_w          <= `ARIANE_CORE204.piton_pc;
                end
            end
    

            assign spc205_thread_id = 2'b00;
            assign spc205_rtl_pc = spc205_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(205*4)]   <= 1'b0;
                  active_thread[(205*4)+1] <= 1'b0;
                  active_thread[(205*4)+2] <= 1'b0;
                  active_thread[(205*4)+3] <= 1'b0;
                  spc205_inst_done         <= 0;
                  spc205_phy_pc_w          <= 0;
                end else begin
                  active_thread[(205*4)]   <= 1'b1;
                  active_thread[(205*4)+1] <= 1'b1;
                  active_thread[(205*4)+2] <= 1'b1;
                  active_thread[(205*4)+3] <= 1'b1;
                  spc205_inst_done         <= `ARIANE_CORE205.piton_pc_vld;
                  spc205_phy_pc_w          <= `ARIANE_CORE205.piton_pc;
                end
            end
    

            assign spc206_thread_id = 2'b00;
            assign spc206_rtl_pc = spc206_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(206*4)]   <= 1'b0;
                  active_thread[(206*4)+1] <= 1'b0;
                  active_thread[(206*4)+2] <= 1'b0;
                  active_thread[(206*4)+3] <= 1'b0;
                  spc206_inst_done         <= 0;
                  spc206_phy_pc_w          <= 0;
                end else begin
                  active_thread[(206*4)]   <= 1'b1;
                  active_thread[(206*4)+1] <= 1'b1;
                  active_thread[(206*4)+2] <= 1'b1;
                  active_thread[(206*4)+3] <= 1'b1;
                  spc206_inst_done         <= `ARIANE_CORE206.piton_pc_vld;
                  spc206_phy_pc_w          <= `ARIANE_CORE206.piton_pc;
                end
            end
    

            assign spc207_thread_id = 2'b00;
            assign spc207_rtl_pc = spc207_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(207*4)]   <= 1'b0;
                  active_thread[(207*4)+1] <= 1'b0;
                  active_thread[(207*4)+2] <= 1'b0;
                  active_thread[(207*4)+3] <= 1'b0;
                  spc207_inst_done         <= 0;
                  spc207_phy_pc_w          <= 0;
                end else begin
                  active_thread[(207*4)]   <= 1'b1;
                  active_thread[(207*4)+1] <= 1'b1;
                  active_thread[(207*4)+2] <= 1'b1;
                  active_thread[(207*4)+3] <= 1'b1;
                  spc207_inst_done         <= `ARIANE_CORE207.piton_pc_vld;
                  spc207_phy_pc_w          <= `ARIANE_CORE207.piton_pc;
                end
            end
    

            assign spc208_thread_id = 2'b00;
            assign spc208_rtl_pc = spc208_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(208*4)]   <= 1'b0;
                  active_thread[(208*4)+1] <= 1'b0;
                  active_thread[(208*4)+2] <= 1'b0;
                  active_thread[(208*4)+3] <= 1'b0;
                  spc208_inst_done         <= 0;
                  spc208_phy_pc_w          <= 0;
                end else begin
                  active_thread[(208*4)]   <= 1'b1;
                  active_thread[(208*4)+1] <= 1'b1;
                  active_thread[(208*4)+2] <= 1'b1;
                  active_thread[(208*4)+3] <= 1'b1;
                  spc208_inst_done         <= `ARIANE_CORE208.piton_pc_vld;
                  spc208_phy_pc_w          <= `ARIANE_CORE208.piton_pc;
                end
            end
    

            assign spc209_thread_id = 2'b00;
            assign spc209_rtl_pc = spc209_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(209*4)]   <= 1'b0;
                  active_thread[(209*4)+1] <= 1'b0;
                  active_thread[(209*4)+2] <= 1'b0;
                  active_thread[(209*4)+3] <= 1'b0;
                  spc209_inst_done         <= 0;
                  spc209_phy_pc_w          <= 0;
                end else begin
                  active_thread[(209*4)]   <= 1'b1;
                  active_thread[(209*4)+1] <= 1'b1;
                  active_thread[(209*4)+2] <= 1'b1;
                  active_thread[(209*4)+3] <= 1'b1;
                  spc209_inst_done         <= `ARIANE_CORE209.piton_pc_vld;
                  spc209_phy_pc_w          <= `ARIANE_CORE209.piton_pc;
                end
            end
    

            assign spc210_thread_id = 2'b00;
            assign spc210_rtl_pc = spc210_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(210*4)]   <= 1'b0;
                  active_thread[(210*4)+1] <= 1'b0;
                  active_thread[(210*4)+2] <= 1'b0;
                  active_thread[(210*4)+3] <= 1'b0;
                  spc210_inst_done         <= 0;
                  spc210_phy_pc_w          <= 0;
                end else begin
                  active_thread[(210*4)]   <= 1'b1;
                  active_thread[(210*4)+1] <= 1'b1;
                  active_thread[(210*4)+2] <= 1'b1;
                  active_thread[(210*4)+3] <= 1'b1;
                  spc210_inst_done         <= `ARIANE_CORE210.piton_pc_vld;
                  spc210_phy_pc_w          <= `ARIANE_CORE210.piton_pc;
                end
            end
    

            assign spc211_thread_id = 2'b00;
            assign spc211_rtl_pc = spc211_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(211*4)]   <= 1'b0;
                  active_thread[(211*4)+1] <= 1'b0;
                  active_thread[(211*4)+2] <= 1'b0;
                  active_thread[(211*4)+3] <= 1'b0;
                  spc211_inst_done         <= 0;
                  spc211_phy_pc_w          <= 0;
                end else begin
                  active_thread[(211*4)]   <= 1'b1;
                  active_thread[(211*4)+1] <= 1'b1;
                  active_thread[(211*4)+2] <= 1'b1;
                  active_thread[(211*4)+3] <= 1'b1;
                  spc211_inst_done         <= `ARIANE_CORE211.piton_pc_vld;
                  spc211_phy_pc_w          <= `ARIANE_CORE211.piton_pc;
                end
            end
    

            assign spc212_thread_id = 2'b00;
            assign spc212_rtl_pc = spc212_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(212*4)]   <= 1'b0;
                  active_thread[(212*4)+1] <= 1'b0;
                  active_thread[(212*4)+2] <= 1'b0;
                  active_thread[(212*4)+3] <= 1'b0;
                  spc212_inst_done         <= 0;
                  spc212_phy_pc_w          <= 0;
                end else begin
                  active_thread[(212*4)]   <= 1'b1;
                  active_thread[(212*4)+1] <= 1'b1;
                  active_thread[(212*4)+2] <= 1'b1;
                  active_thread[(212*4)+3] <= 1'b1;
                  spc212_inst_done         <= `ARIANE_CORE212.piton_pc_vld;
                  spc212_phy_pc_w          <= `ARIANE_CORE212.piton_pc;
                end
            end
    

            assign spc213_thread_id = 2'b00;
            assign spc213_rtl_pc = spc213_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(213*4)]   <= 1'b0;
                  active_thread[(213*4)+1] <= 1'b0;
                  active_thread[(213*4)+2] <= 1'b0;
                  active_thread[(213*4)+3] <= 1'b0;
                  spc213_inst_done         <= 0;
                  spc213_phy_pc_w          <= 0;
                end else begin
                  active_thread[(213*4)]   <= 1'b1;
                  active_thread[(213*4)+1] <= 1'b1;
                  active_thread[(213*4)+2] <= 1'b1;
                  active_thread[(213*4)+3] <= 1'b1;
                  spc213_inst_done         <= `ARIANE_CORE213.piton_pc_vld;
                  spc213_phy_pc_w          <= `ARIANE_CORE213.piton_pc;
                end
            end
    

            assign spc214_thread_id = 2'b00;
            assign spc214_rtl_pc = spc214_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(214*4)]   <= 1'b0;
                  active_thread[(214*4)+1] <= 1'b0;
                  active_thread[(214*4)+2] <= 1'b0;
                  active_thread[(214*4)+3] <= 1'b0;
                  spc214_inst_done         <= 0;
                  spc214_phy_pc_w          <= 0;
                end else begin
                  active_thread[(214*4)]   <= 1'b1;
                  active_thread[(214*4)+1] <= 1'b1;
                  active_thread[(214*4)+2] <= 1'b1;
                  active_thread[(214*4)+3] <= 1'b1;
                  spc214_inst_done         <= `ARIANE_CORE214.piton_pc_vld;
                  spc214_phy_pc_w          <= `ARIANE_CORE214.piton_pc;
                end
            end
    

            assign spc215_thread_id = 2'b00;
            assign spc215_rtl_pc = spc215_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(215*4)]   <= 1'b0;
                  active_thread[(215*4)+1] <= 1'b0;
                  active_thread[(215*4)+2] <= 1'b0;
                  active_thread[(215*4)+3] <= 1'b0;
                  spc215_inst_done         <= 0;
                  spc215_phy_pc_w          <= 0;
                end else begin
                  active_thread[(215*4)]   <= 1'b1;
                  active_thread[(215*4)+1] <= 1'b1;
                  active_thread[(215*4)+2] <= 1'b1;
                  active_thread[(215*4)+3] <= 1'b1;
                  spc215_inst_done         <= `ARIANE_CORE215.piton_pc_vld;
                  spc215_phy_pc_w          <= `ARIANE_CORE215.piton_pc;
                end
            end
    

            assign spc216_thread_id = 2'b00;
            assign spc216_rtl_pc = spc216_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(216*4)]   <= 1'b0;
                  active_thread[(216*4)+1] <= 1'b0;
                  active_thread[(216*4)+2] <= 1'b0;
                  active_thread[(216*4)+3] <= 1'b0;
                  spc216_inst_done         <= 0;
                  spc216_phy_pc_w          <= 0;
                end else begin
                  active_thread[(216*4)]   <= 1'b1;
                  active_thread[(216*4)+1] <= 1'b1;
                  active_thread[(216*4)+2] <= 1'b1;
                  active_thread[(216*4)+3] <= 1'b1;
                  spc216_inst_done         <= `ARIANE_CORE216.piton_pc_vld;
                  spc216_phy_pc_w          <= `ARIANE_CORE216.piton_pc;
                end
            end
    

            assign spc217_thread_id = 2'b00;
            assign spc217_rtl_pc = spc217_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(217*4)]   <= 1'b0;
                  active_thread[(217*4)+1] <= 1'b0;
                  active_thread[(217*4)+2] <= 1'b0;
                  active_thread[(217*4)+3] <= 1'b0;
                  spc217_inst_done         <= 0;
                  spc217_phy_pc_w          <= 0;
                end else begin
                  active_thread[(217*4)]   <= 1'b1;
                  active_thread[(217*4)+1] <= 1'b1;
                  active_thread[(217*4)+2] <= 1'b1;
                  active_thread[(217*4)+3] <= 1'b1;
                  spc217_inst_done         <= `ARIANE_CORE217.piton_pc_vld;
                  spc217_phy_pc_w          <= `ARIANE_CORE217.piton_pc;
                end
            end
    

            assign spc218_thread_id = 2'b00;
            assign spc218_rtl_pc = spc218_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(218*4)]   <= 1'b0;
                  active_thread[(218*4)+1] <= 1'b0;
                  active_thread[(218*4)+2] <= 1'b0;
                  active_thread[(218*4)+3] <= 1'b0;
                  spc218_inst_done         <= 0;
                  spc218_phy_pc_w          <= 0;
                end else begin
                  active_thread[(218*4)]   <= 1'b1;
                  active_thread[(218*4)+1] <= 1'b1;
                  active_thread[(218*4)+2] <= 1'b1;
                  active_thread[(218*4)+3] <= 1'b1;
                  spc218_inst_done         <= `ARIANE_CORE218.piton_pc_vld;
                  spc218_phy_pc_w          <= `ARIANE_CORE218.piton_pc;
                end
            end
    

            assign spc219_thread_id = 2'b00;
            assign spc219_rtl_pc = spc219_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(219*4)]   <= 1'b0;
                  active_thread[(219*4)+1] <= 1'b0;
                  active_thread[(219*4)+2] <= 1'b0;
                  active_thread[(219*4)+3] <= 1'b0;
                  spc219_inst_done         <= 0;
                  spc219_phy_pc_w          <= 0;
                end else begin
                  active_thread[(219*4)]   <= 1'b1;
                  active_thread[(219*4)+1] <= 1'b1;
                  active_thread[(219*4)+2] <= 1'b1;
                  active_thread[(219*4)+3] <= 1'b1;
                  spc219_inst_done         <= `ARIANE_CORE219.piton_pc_vld;
                  spc219_phy_pc_w          <= `ARIANE_CORE219.piton_pc;
                end
            end
    

            assign spc220_thread_id = 2'b00;
            assign spc220_rtl_pc = spc220_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(220*4)]   <= 1'b0;
                  active_thread[(220*4)+1] <= 1'b0;
                  active_thread[(220*4)+2] <= 1'b0;
                  active_thread[(220*4)+3] <= 1'b0;
                  spc220_inst_done         <= 0;
                  spc220_phy_pc_w          <= 0;
                end else begin
                  active_thread[(220*4)]   <= 1'b1;
                  active_thread[(220*4)+1] <= 1'b1;
                  active_thread[(220*4)+2] <= 1'b1;
                  active_thread[(220*4)+3] <= 1'b1;
                  spc220_inst_done         <= `ARIANE_CORE220.piton_pc_vld;
                  spc220_phy_pc_w          <= `ARIANE_CORE220.piton_pc;
                end
            end
    

            assign spc221_thread_id = 2'b00;
            assign spc221_rtl_pc = spc221_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(221*4)]   <= 1'b0;
                  active_thread[(221*4)+1] <= 1'b0;
                  active_thread[(221*4)+2] <= 1'b0;
                  active_thread[(221*4)+3] <= 1'b0;
                  spc221_inst_done         <= 0;
                  spc221_phy_pc_w          <= 0;
                end else begin
                  active_thread[(221*4)]   <= 1'b1;
                  active_thread[(221*4)+1] <= 1'b1;
                  active_thread[(221*4)+2] <= 1'b1;
                  active_thread[(221*4)+3] <= 1'b1;
                  spc221_inst_done         <= `ARIANE_CORE221.piton_pc_vld;
                  spc221_phy_pc_w          <= `ARIANE_CORE221.piton_pc;
                end
            end
    

            assign spc222_thread_id = 2'b00;
            assign spc222_rtl_pc = spc222_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(222*4)]   <= 1'b0;
                  active_thread[(222*4)+1] <= 1'b0;
                  active_thread[(222*4)+2] <= 1'b0;
                  active_thread[(222*4)+3] <= 1'b0;
                  spc222_inst_done         <= 0;
                  spc222_phy_pc_w          <= 0;
                end else begin
                  active_thread[(222*4)]   <= 1'b1;
                  active_thread[(222*4)+1] <= 1'b1;
                  active_thread[(222*4)+2] <= 1'b1;
                  active_thread[(222*4)+3] <= 1'b1;
                  spc222_inst_done         <= `ARIANE_CORE222.piton_pc_vld;
                  spc222_phy_pc_w          <= `ARIANE_CORE222.piton_pc;
                end
            end
    

            assign spc223_thread_id = 2'b00;
            assign spc223_rtl_pc = spc223_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(223*4)]   <= 1'b0;
                  active_thread[(223*4)+1] <= 1'b0;
                  active_thread[(223*4)+2] <= 1'b0;
                  active_thread[(223*4)+3] <= 1'b0;
                  spc223_inst_done         <= 0;
                  spc223_phy_pc_w          <= 0;
                end else begin
                  active_thread[(223*4)]   <= 1'b1;
                  active_thread[(223*4)+1] <= 1'b1;
                  active_thread[(223*4)+2] <= 1'b1;
                  active_thread[(223*4)+3] <= 1'b1;
                  spc223_inst_done         <= `ARIANE_CORE223.piton_pc_vld;
                  spc223_phy_pc_w          <= `ARIANE_CORE223.piton_pc;
                end
            end
    

            assign spc224_thread_id = 2'b00;
            assign spc224_rtl_pc = spc224_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(224*4)]   <= 1'b0;
                  active_thread[(224*4)+1] <= 1'b0;
                  active_thread[(224*4)+2] <= 1'b0;
                  active_thread[(224*4)+3] <= 1'b0;
                  spc224_inst_done         <= 0;
                  spc224_phy_pc_w          <= 0;
                end else begin
                  active_thread[(224*4)]   <= 1'b1;
                  active_thread[(224*4)+1] <= 1'b1;
                  active_thread[(224*4)+2] <= 1'b1;
                  active_thread[(224*4)+3] <= 1'b1;
                  spc224_inst_done         <= `ARIANE_CORE224.piton_pc_vld;
                  spc224_phy_pc_w          <= `ARIANE_CORE224.piton_pc;
                end
            end
    

            assign spc225_thread_id = 2'b00;
            assign spc225_rtl_pc = spc225_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(225*4)]   <= 1'b0;
                  active_thread[(225*4)+1] <= 1'b0;
                  active_thread[(225*4)+2] <= 1'b0;
                  active_thread[(225*4)+3] <= 1'b0;
                  spc225_inst_done         <= 0;
                  spc225_phy_pc_w          <= 0;
                end else begin
                  active_thread[(225*4)]   <= 1'b1;
                  active_thread[(225*4)+1] <= 1'b1;
                  active_thread[(225*4)+2] <= 1'b1;
                  active_thread[(225*4)+3] <= 1'b1;
                  spc225_inst_done         <= `ARIANE_CORE225.piton_pc_vld;
                  spc225_phy_pc_w          <= `ARIANE_CORE225.piton_pc;
                end
            end
    

            assign spc226_thread_id = 2'b00;
            assign spc226_rtl_pc = spc226_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(226*4)]   <= 1'b0;
                  active_thread[(226*4)+1] <= 1'b0;
                  active_thread[(226*4)+2] <= 1'b0;
                  active_thread[(226*4)+3] <= 1'b0;
                  spc226_inst_done         <= 0;
                  spc226_phy_pc_w          <= 0;
                end else begin
                  active_thread[(226*4)]   <= 1'b1;
                  active_thread[(226*4)+1] <= 1'b1;
                  active_thread[(226*4)+2] <= 1'b1;
                  active_thread[(226*4)+3] <= 1'b1;
                  spc226_inst_done         <= `ARIANE_CORE226.piton_pc_vld;
                  spc226_phy_pc_w          <= `ARIANE_CORE226.piton_pc;
                end
            end
    

            assign spc227_thread_id = 2'b00;
            assign spc227_rtl_pc = spc227_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(227*4)]   <= 1'b0;
                  active_thread[(227*4)+1] <= 1'b0;
                  active_thread[(227*4)+2] <= 1'b0;
                  active_thread[(227*4)+3] <= 1'b0;
                  spc227_inst_done         <= 0;
                  spc227_phy_pc_w          <= 0;
                end else begin
                  active_thread[(227*4)]   <= 1'b1;
                  active_thread[(227*4)+1] <= 1'b1;
                  active_thread[(227*4)+2] <= 1'b1;
                  active_thread[(227*4)+3] <= 1'b1;
                  spc227_inst_done         <= `ARIANE_CORE227.piton_pc_vld;
                  spc227_phy_pc_w          <= `ARIANE_CORE227.piton_pc;
                end
            end
    

            assign spc228_thread_id = 2'b00;
            assign spc228_rtl_pc = spc228_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(228*4)]   <= 1'b0;
                  active_thread[(228*4)+1] <= 1'b0;
                  active_thread[(228*4)+2] <= 1'b0;
                  active_thread[(228*4)+3] <= 1'b0;
                  spc228_inst_done         <= 0;
                  spc228_phy_pc_w          <= 0;
                end else begin
                  active_thread[(228*4)]   <= 1'b1;
                  active_thread[(228*4)+1] <= 1'b1;
                  active_thread[(228*4)+2] <= 1'b1;
                  active_thread[(228*4)+3] <= 1'b1;
                  spc228_inst_done         <= `ARIANE_CORE228.piton_pc_vld;
                  spc228_phy_pc_w          <= `ARIANE_CORE228.piton_pc;
                end
            end
    

            assign spc229_thread_id = 2'b00;
            assign spc229_rtl_pc = spc229_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(229*4)]   <= 1'b0;
                  active_thread[(229*4)+1] <= 1'b0;
                  active_thread[(229*4)+2] <= 1'b0;
                  active_thread[(229*4)+3] <= 1'b0;
                  spc229_inst_done         <= 0;
                  spc229_phy_pc_w          <= 0;
                end else begin
                  active_thread[(229*4)]   <= 1'b1;
                  active_thread[(229*4)+1] <= 1'b1;
                  active_thread[(229*4)+2] <= 1'b1;
                  active_thread[(229*4)+3] <= 1'b1;
                  spc229_inst_done         <= `ARIANE_CORE229.piton_pc_vld;
                  spc229_phy_pc_w          <= `ARIANE_CORE229.piton_pc;
                end
            end
    

            assign spc230_thread_id = 2'b00;
            assign spc230_rtl_pc = spc230_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(230*4)]   <= 1'b0;
                  active_thread[(230*4)+1] <= 1'b0;
                  active_thread[(230*4)+2] <= 1'b0;
                  active_thread[(230*4)+3] <= 1'b0;
                  spc230_inst_done         <= 0;
                  spc230_phy_pc_w          <= 0;
                end else begin
                  active_thread[(230*4)]   <= 1'b1;
                  active_thread[(230*4)+1] <= 1'b1;
                  active_thread[(230*4)+2] <= 1'b1;
                  active_thread[(230*4)+3] <= 1'b1;
                  spc230_inst_done         <= `ARIANE_CORE230.piton_pc_vld;
                  spc230_phy_pc_w          <= `ARIANE_CORE230.piton_pc;
                end
            end
    

            assign spc231_thread_id = 2'b00;
            assign spc231_rtl_pc = spc231_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(231*4)]   <= 1'b0;
                  active_thread[(231*4)+1] <= 1'b0;
                  active_thread[(231*4)+2] <= 1'b0;
                  active_thread[(231*4)+3] <= 1'b0;
                  spc231_inst_done         <= 0;
                  spc231_phy_pc_w          <= 0;
                end else begin
                  active_thread[(231*4)]   <= 1'b1;
                  active_thread[(231*4)+1] <= 1'b1;
                  active_thread[(231*4)+2] <= 1'b1;
                  active_thread[(231*4)+3] <= 1'b1;
                  spc231_inst_done         <= `ARIANE_CORE231.piton_pc_vld;
                  spc231_phy_pc_w          <= `ARIANE_CORE231.piton_pc;
                end
            end
    

            assign spc232_thread_id = 2'b00;
            assign spc232_rtl_pc = spc232_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(232*4)]   <= 1'b0;
                  active_thread[(232*4)+1] <= 1'b0;
                  active_thread[(232*4)+2] <= 1'b0;
                  active_thread[(232*4)+3] <= 1'b0;
                  spc232_inst_done         <= 0;
                  spc232_phy_pc_w          <= 0;
                end else begin
                  active_thread[(232*4)]   <= 1'b1;
                  active_thread[(232*4)+1] <= 1'b1;
                  active_thread[(232*4)+2] <= 1'b1;
                  active_thread[(232*4)+3] <= 1'b1;
                  spc232_inst_done         <= `ARIANE_CORE232.piton_pc_vld;
                  spc232_phy_pc_w          <= `ARIANE_CORE232.piton_pc;
                end
            end
    

            assign spc233_thread_id = 2'b00;
            assign spc233_rtl_pc = spc233_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(233*4)]   <= 1'b0;
                  active_thread[(233*4)+1] <= 1'b0;
                  active_thread[(233*4)+2] <= 1'b0;
                  active_thread[(233*4)+3] <= 1'b0;
                  spc233_inst_done         <= 0;
                  spc233_phy_pc_w          <= 0;
                end else begin
                  active_thread[(233*4)]   <= 1'b1;
                  active_thread[(233*4)+1] <= 1'b1;
                  active_thread[(233*4)+2] <= 1'b1;
                  active_thread[(233*4)+3] <= 1'b1;
                  spc233_inst_done         <= `ARIANE_CORE233.piton_pc_vld;
                  spc233_phy_pc_w          <= `ARIANE_CORE233.piton_pc;
                end
            end
    

            assign spc234_thread_id = 2'b00;
            assign spc234_rtl_pc = spc234_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(234*4)]   <= 1'b0;
                  active_thread[(234*4)+1] <= 1'b0;
                  active_thread[(234*4)+2] <= 1'b0;
                  active_thread[(234*4)+3] <= 1'b0;
                  spc234_inst_done         <= 0;
                  spc234_phy_pc_w          <= 0;
                end else begin
                  active_thread[(234*4)]   <= 1'b1;
                  active_thread[(234*4)+1] <= 1'b1;
                  active_thread[(234*4)+2] <= 1'b1;
                  active_thread[(234*4)+3] <= 1'b1;
                  spc234_inst_done         <= `ARIANE_CORE234.piton_pc_vld;
                  spc234_phy_pc_w          <= `ARIANE_CORE234.piton_pc;
                end
            end
    

            assign spc235_thread_id = 2'b00;
            assign spc235_rtl_pc = spc235_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(235*4)]   <= 1'b0;
                  active_thread[(235*4)+1] <= 1'b0;
                  active_thread[(235*4)+2] <= 1'b0;
                  active_thread[(235*4)+3] <= 1'b0;
                  spc235_inst_done         <= 0;
                  spc235_phy_pc_w          <= 0;
                end else begin
                  active_thread[(235*4)]   <= 1'b1;
                  active_thread[(235*4)+1] <= 1'b1;
                  active_thread[(235*4)+2] <= 1'b1;
                  active_thread[(235*4)+3] <= 1'b1;
                  spc235_inst_done         <= `ARIANE_CORE235.piton_pc_vld;
                  spc235_phy_pc_w          <= `ARIANE_CORE235.piton_pc;
                end
            end
    

            assign spc236_thread_id = 2'b00;
            assign spc236_rtl_pc = spc236_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(236*4)]   <= 1'b0;
                  active_thread[(236*4)+1] <= 1'b0;
                  active_thread[(236*4)+2] <= 1'b0;
                  active_thread[(236*4)+3] <= 1'b0;
                  spc236_inst_done         <= 0;
                  spc236_phy_pc_w          <= 0;
                end else begin
                  active_thread[(236*4)]   <= 1'b1;
                  active_thread[(236*4)+1] <= 1'b1;
                  active_thread[(236*4)+2] <= 1'b1;
                  active_thread[(236*4)+3] <= 1'b1;
                  spc236_inst_done         <= `ARIANE_CORE236.piton_pc_vld;
                  spc236_phy_pc_w          <= `ARIANE_CORE236.piton_pc;
                end
            end
    

            assign spc237_thread_id = 2'b00;
            assign spc237_rtl_pc = spc237_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(237*4)]   <= 1'b0;
                  active_thread[(237*4)+1] <= 1'b0;
                  active_thread[(237*4)+2] <= 1'b0;
                  active_thread[(237*4)+3] <= 1'b0;
                  spc237_inst_done         <= 0;
                  spc237_phy_pc_w          <= 0;
                end else begin
                  active_thread[(237*4)]   <= 1'b1;
                  active_thread[(237*4)+1] <= 1'b1;
                  active_thread[(237*4)+2] <= 1'b1;
                  active_thread[(237*4)+3] <= 1'b1;
                  spc237_inst_done         <= `ARIANE_CORE237.piton_pc_vld;
                  spc237_phy_pc_w          <= `ARIANE_CORE237.piton_pc;
                end
            end
    

            assign spc238_thread_id = 2'b00;
            assign spc238_rtl_pc = spc238_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(238*4)]   <= 1'b0;
                  active_thread[(238*4)+1] <= 1'b0;
                  active_thread[(238*4)+2] <= 1'b0;
                  active_thread[(238*4)+3] <= 1'b0;
                  spc238_inst_done         <= 0;
                  spc238_phy_pc_w          <= 0;
                end else begin
                  active_thread[(238*4)]   <= 1'b1;
                  active_thread[(238*4)+1] <= 1'b1;
                  active_thread[(238*4)+2] <= 1'b1;
                  active_thread[(238*4)+3] <= 1'b1;
                  spc238_inst_done         <= `ARIANE_CORE238.piton_pc_vld;
                  spc238_phy_pc_w          <= `ARIANE_CORE238.piton_pc;
                end
            end
    

            assign spc239_thread_id = 2'b00;
            assign spc239_rtl_pc = spc239_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(239*4)]   <= 1'b0;
                  active_thread[(239*4)+1] <= 1'b0;
                  active_thread[(239*4)+2] <= 1'b0;
                  active_thread[(239*4)+3] <= 1'b0;
                  spc239_inst_done         <= 0;
                  spc239_phy_pc_w          <= 0;
                end else begin
                  active_thread[(239*4)]   <= 1'b1;
                  active_thread[(239*4)+1] <= 1'b1;
                  active_thread[(239*4)+2] <= 1'b1;
                  active_thread[(239*4)+3] <= 1'b1;
                  spc239_inst_done         <= `ARIANE_CORE239.piton_pc_vld;
                  spc239_phy_pc_w          <= `ARIANE_CORE239.piton_pc;
                end
            end
    

            assign spc240_thread_id = 2'b00;
            assign spc240_rtl_pc = spc240_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(240*4)]   <= 1'b0;
                  active_thread[(240*4)+1] <= 1'b0;
                  active_thread[(240*4)+2] <= 1'b0;
                  active_thread[(240*4)+3] <= 1'b0;
                  spc240_inst_done         <= 0;
                  spc240_phy_pc_w          <= 0;
                end else begin
                  active_thread[(240*4)]   <= 1'b1;
                  active_thread[(240*4)+1] <= 1'b1;
                  active_thread[(240*4)+2] <= 1'b1;
                  active_thread[(240*4)+3] <= 1'b1;
                  spc240_inst_done         <= `ARIANE_CORE240.piton_pc_vld;
                  spc240_phy_pc_w          <= `ARIANE_CORE240.piton_pc;
                end
            end
    

            assign spc241_thread_id = 2'b00;
            assign spc241_rtl_pc = spc241_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(241*4)]   <= 1'b0;
                  active_thread[(241*4)+1] <= 1'b0;
                  active_thread[(241*4)+2] <= 1'b0;
                  active_thread[(241*4)+3] <= 1'b0;
                  spc241_inst_done         <= 0;
                  spc241_phy_pc_w          <= 0;
                end else begin
                  active_thread[(241*4)]   <= 1'b1;
                  active_thread[(241*4)+1] <= 1'b1;
                  active_thread[(241*4)+2] <= 1'b1;
                  active_thread[(241*4)+3] <= 1'b1;
                  spc241_inst_done         <= `ARIANE_CORE241.piton_pc_vld;
                  spc241_phy_pc_w          <= `ARIANE_CORE241.piton_pc;
                end
            end
    

            assign spc242_thread_id = 2'b00;
            assign spc242_rtl_pc = spc242_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(242*4)]   <= 1'b0;
                  active_thread[(242*4)+1] <= 1'b0;
                  active_thread[(242*4)+2] <= 1'b0;
                  active_thread[(242*4)+3] <= 1'b0;
                  spc242_inst_done         <= 0;
                  spc242_phy_pc_w          <= 0;
                end else begin
                  active_thread[(242*4)]   <= 1'b1;
                  active_thread[(242*4)+1] <= 1'b1;
                  active_thread[(242*4)+2] <= 1'b1;
                  active_thread[(242*4)+3] <= 1'b1;
                  spc242_inst_done         <= `ARIANE_CORE242.piton_pc_vld;
                  spc242_phy_pc_w          <= `ARIANE_CORE242.piton_pc;
                end
            end
    

            assign spc243_thread_id = 2'b00;
            assign spc243_rtl_pc = spc243_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(243*4)]   <= 1'b0;
                  active_thread[(243*4)+1] <= 1'b0;
                  active_thread[(243*4)+2] <= 1'b0;
                  active_thread[(243*4)+3] <= 1'b0;
                  spc243_inst_done         <= 0;
                  spc243_phy_pc_w          <= 0;
                end else begin
                  active_thread[(243*4)]   <= 1'b1;
                  active_thread[(243*4)+1] <= 1'b1;
                  active_thread[(243*4)+2] <= 1'b1;
                  active_thread[(243*4)+3] <= 1'b1;
                  spc243_inst_done         <= `ARIANE_CORE243.piton_pc_vld;
                  spc243_phy_pc_w          <= `ARIANE_CORE243.piton_pc;
                end
            end
    

            assign spc244_thread_id = 2'b00;
            assign spc244_rtl_pc = spc244_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(244*4)]   <= 1'b0;
                  active_thread[(244*4)+1] <= 1'b0;
                  active_thread[(244*4)+2] <= 1'b0;
                  active_thread[(244*4)+3] <= 1'b0;
                  spc244_inst_done         <= 0;
                  spc244_phy_pc_w          <= 0;
                end else begin
                  active_thread[(244*4)]   <= 1'b1;
                  active_thread[(244*4)+1] <= 1'b1;
                  active_thread[(244*4)+2] <= 1'b1;
                  active_thread[(244*4)+3] <= 1'b1;
                  spc244_inst_done         <= `ARIANE_CORE244.piton_pc_vld;
                  spc244_phy_pc_w          <= `ARIANE_CORE244.piton_pc;
                end
            end
    

            assign spc245_thread_id = 2'b00;
            assign spc245_rtl_pc = spc245_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(245*4)]   <= 1'b0;
                  active_thread[(245*4)+1] <= 1'b0;
                  active_thread[(245*4)+2] <= 1'b0;
                  active_thread[(245*4)+3] <= 1'b0;
                  spc245_inst_done         <= 0;
                  spc245_phy_pc_w          <= 0;
                end else begin
                  active_thread[(245*4)]   <= 1'b1;
                  active_thread[(245*4)+1] <= 1'b1;
                  active_thread[(245*4)+2] <= 1'b1;
                  active_thread[(245*4)+3] <= 1'b1;
                  spc245_inst_done         <= `ARIANE_CORE245.piton_pc_vld;
                  spc245_phy_pc_w          <= `ARIANE_CORE245.piton_pc;
                end
            end
    

            assign spc246_thread_id = 2'b00;
            assign spc246_rtl_pc = spc246_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(246*4)]   <= 1'b0;
                  active_thread[(246*4)+1] <= 1'b0;
                  active_thread[(246*4)+2] <= 1'b0;
                  active_thread[(246*4)+3] <= 1'b0;
                  spc246_inst_done         <= 0;
                  spc246_phy_pc_w          <= 0;
                end else begin
                  active_thread[(246*4)]   <= 1'b1;
                  active_thread[(246*4)+1] <= 1'b1;
                  active_thread[(246*4)+2] <= 1'b1;
                  active_thread[(246*4)+3] <= 1'b1;
                  spc246_inst_done         <= `ARIANE_CORE246.piton_pc_vld;
                  spc246_phy_pc_w          <= `ARIANE_CORE246.piton_pc;
                end
            end
    

            assign spc247_thread_id = 2'b00;
            assign spc247_rtl_pc = spc247_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(247*4)]   <= 1'b0;
                  active_thread[(247*4)+1] <= 1'b0;
                  active_thread[(247*4)+2] <= 1'b0;
                  active_thread[(247*4)+3] <= 1'b0;
                  spc247_inst_done         <= 0;
                  spc247_phy_pc_w          <= 0;
                end else begin
                  active_thread[(247*4)]   <= 1'b1;
                  active_thread[(247*4)+1] <= 1'b1;
                  active_thread[(247*4)+2] <= 1'b1;
                  active_thread[(247*4)+3] <= 1'b1;
                  spc247_inst_done         <= `ARIANE_CORE247.piton_pc_vld;
                  spc247_phy_pc_w          <= `ARIANE_CORE247.piton_pc;
                end
            end
    

            assign spc248_thread_id = 2'b00;
            assign spc248_rtl_pc = spc248_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(248*4)]   <= 1'b0;
                  active_thread[(248*4)+1] <= 1'b0;
                  active_thread[(248*4)+2] <= 1'b0;
                  active_thread[(248*4)+3] <= 1'b0;
                  spc248_inst_done         <= 0;
                  spc248_phy_pc_w          <= 0;
                end else begin
                  active_thread[(248*4)]   <= 1'b1;
                  active_thread[(248*4)+1] <= 1'b1;
                  active_thread[(248*4)+2] <= 1'b1;
                  active_thread[(248*4)+3] <= 1'b1;
                  spc248_inst_done         <= `ARIANE_CORE248.piton_pc_vld;
                  spc248_phy_pc_w          <= `ARIANE_CORE248.piton_pc;
                end
            end
    

            assign spc249_thread_id = 2'b00;
            assign spc249_rtl_pc = spc249_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(249*4)]   <= 1'b0;
                  active_thread[(249*4)+1] <= 1'b0;
                  active_thread[(249*4)+2] <= 1'b0;
                  active_thread[(249*4)+3] <= 1'b0;
                  spc249_inst_done         <= 0;
                  spc249_phy_pc_w          <= 0;
                end else begin
                  active_thread[(249*4)]   <= 1'b1;
                  active_thread[(249*4)+1] <= 1'b1;
                  active_thread[(249*4)+2] <= 1'b1;
                  active_thread[(249*4)+3] <= 1'b1;
                  spc249_inst_done         <= `ARIANE_CORE249.piton_pc_vld;
                  spc249_phy_pc_w          <= `ARIANE_CORE249.piton_pc;
                end
            end
    

            assign spc250_thread_id = 2'b00;
            assign spc250_rtl_pc = spc250_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(250*4)]   <= 1'b0;
                  active_thread[(250*4)+1] <= 1'b0;
                  active_thread[(250*4)+2] <= 1'b0;
                  active_thread[(250*4)+3] <= 1'b0;
                  spc250_inst_done         <= 0;
                  spc250_phy_pc_w          <= 0;
                end else begin
                  active_thread[(250*4)]   <= 1'b1;
                  active_thread[(250*4)+1] <= 1'b1;
                  active_thread[(250*4)+2] <= 1'b1;
                  active_thread[(250*4)+3] <= 1'b1;
                  spc250_inst_done         <= `ARIANE_CORE250.piton_pc_vld;
                  spc250_phy_pc_w          <= `ARIANE_CORE250.piton_pc;
                end
            end
    

            assign spc251_thread_id = 2'b00;
            assign spc251_rtl_pc = spc251_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(251*4)]   <= 1'b0;
                  active_thread[(251*4)+1] <= 1'b0;
                  active_thread[(251*4)+2] <= 1'b0;
                  active_thread[(251*4)+3] <= 1'b0;
                  spc251_inst_done         <= 0;
                  spc251_phy_pc_w          <= 0;
                end else begin
                  active_thread[(251*4)]   <= 1'b1;
                  active_thread[(251*4)+1] <= 1'b1;
                  active_thread[(251*4)+2] <= 1'b1;
                  active_thread[(251*4)+3] <= 1'b1;
                  spc251_inst_done         <= `ARIANE_CORE251.piton_pc_vld;
                  spc251_phy_pc_w          <= `ARIANE_CORE251.piton_pc;
                end
            end
    

            assign spc252_thread_id = 2'b00;
            assign spc252_rtl_pc = spc252_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(252*4)]   <= 1'b0;
                  active_thread[(252*4)+1] <= 1'b0;
                  active_thread[(252*4)+2] <= 1'b0;
                  active_thread[(252*4)+3] <= 1'b0;
                  spc252_inst_done         <= 0;
                  spc252_phy_pc_w          <= 0;
                end else begin
                  active_thread[(252*4)]   <= 1'b1;
                  active_thread[(252*4)+1] <= 1'b1;
                  active_thread[(252*4)+2] <= 1'b1;
                  active_thread[(252*4)+3] <= 1'b1;
                  spc252_inst_done         <= `ARIANE_CORE252.piton_pc_vld;
                  spc252_phy_pc_w          <= `ARIANE_CORE252.piton_pc;
                end
            end
    

            assign spc253_thread_id = 2'b00;
            assign spc253_rtl_pc = spc253_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(253*4)]   <= 1'b0;
                  active_thread[(253*4)+1] <= 1'b0;
                  active_thread[(253*4)+2] <= 1'b0;
                  active_thread[(253*4)+3] <= 1'b0;
                  spc253_inst_done         <= 0;
                  spc253_phy_pc_w          <= 0;
                end else begin
                  active_thread[(253*4)]   <= 1'b1;
                  active_thread[(253*4)+1] <= 1'b1;
                  active_thread[(253*4)+2] <= 1'b1;
                  active_thread[(253*4)+3] <= 1'b1;
                  spc253_inst_done         <= `ARIANE_CORE253.piton_pc_vld;
                  spc253_phy_pc_w          <= `ARIANE_CORE253.piton_pc;
                end
            end
    

            assign spc254_thread_id = 2'b00;
            assign spc254_rtl_pc = spc254_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(254*4)]   <= 1'b0;
                  active_thread[(254*4)+1] <= 1'b0;
                  active_thread[(254*4)+2] <= 1'b0;
                  active_thread[(254*4)+3] <= 1'b0;
                  spc254_inst_done         <= 0;
                  spc254_phy_pc_w          <= 0;
                end else begin
                  active_thread[(254*4)]   <= 1'b1;
                  active_thread[(254*4)+1] <= 1'b1;
                  active_thread[(254*4)+2] <= 1'b1;
                  active_thread[(254*4)+3] <= 1'b1;
                  spc254_inst_done         <= `ARIANE_CORE254.piton_pc_vld;
                  spc254_phy_pc_w          <= `ARIANE_CORE254.piton_pc;
                end
            end
    

            assign spc255_thread_id = 2'b00;
            assign spc255_rtl_pc = spc255_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(255*4)]   <= 1'b0;
                  active_thread[(255*4)+1] <= 1'b0;
                  active_thread[(255*4)+2] <= 1'b0;
                  active_thread[(255*4)+3] <= 1'b0;
                  spc255_inst_done         <= 0;
                  spc255_phy_pc_w          <= 0;
                end else begin
                  active_thread[(255*4)]   <= 1'b1;
                  active_thread[(255*4)+1] <= 1'b1;
                  active_thread[(255*4)+2] <= 1'b1;
                  active_thread[(255*4)+3] <= 1'b1;
                  spc255_inst_done         <= `ARIANE_CORE255.piton_pc_vld;
                  spc255_phy_pc_w          <= `ARIANE_CORE255.piton_pc;
                end
            end
    

            assign spc256_thread_id = 2'b00;
            assign spc256_rtl_pc = spc256_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(256*4)]   <= 1'b0;
                  active_thread[(256*4)+1] <= 1'b0;
                  active_thread[(256*4)+2] <= 1'b0;
                  active_thread[(256*4)+3] <= 1'b0;
                  spc256_inst_done         <= 0;
                  spc256_phy_pc_w          <= 0;
                end else begin
                  active_thread[(256*4)]   <= 1'b1;
                  active_thread[(256*4)+1] <= 1'b1;
                  active_thread[(256*4)+2] <= 1'b1;
                  active_thread[(256*4)+3] <= 1'b1;
                  spc256_inst_done         <= `ARIANE_CORE256.piton_pc_vld;
                  spc256_phy_pc_w          <= `ARIANE_CORE256.piton_pc;
                end
            end
    

            assign spc257_thread_id = 2'b00;
            assign spc257_rtl_pc = spc257_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(257*4)]   <= 1'b0;
                  active_thread[(257*4)+1] <= 1'b0;
                  active_thread[(257*4)+2] <= 1'b0;
                  active_thread[(257*4)+3] <= 1'b0;
                  spc257_inst_done         <= 0;
                  spc257_phy_pc_w          <= 0;
                end else begin
                  active_thread[(257*4)]   <= 1'b1;
                  active_thread[(257*4)+1] <= 1'b1;
                  active_thread[(257*4)+2] <= 1'b1;
                  active_thread[(257*4)+3] <= 1'b1;
                  spc257_inst_done         <= `ARIANE_CORE257.piton_pc_vld;
                  spc257_phy_pc_w          <= `ARIANE_CORE257.piton_pc;
                end
            end
    

            assign spc258_thread_id = 2'b00;
            assign spc258_rtl_pc = spc258_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(258*4)]   <= 1'b0;
                  active_thread[(258*4)+1] <= 1'b0;
                  active_thread[(258*4)+2] <= 1'b0;
                  active_thread[(258*4)+3] <= 1'b0;
                  spc258_inst_done         <= 0;
                  spc258_phy_pc_w          <= 0;
                end else begin
                  active_thread[(258*4)]   <= 1'b1;
                  active_thread[(258*4)+1] <= 1'b1;
                  active_thread[(258*4)+2] <= 1'b1;
                  active_thread[(258*4)+3] <= 1'b1;
                  spc258_inst_done         <= `ARIANE_CORE258.piton_pc_vld;
                  spc258_phy_pc_w          <= `ARIANE_CORE258.piton_pc;
                end
            end
    

            assign spc259_thread_id = 2'b00;
            assign spc259_rtl_pc = spc259_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(259*4)]   <= 1'b0;
                  active_thread[(259*4)+1] <= 1'b0;
                  active_thread[(259*4)+2] <= 1'b0;
                  active_thread[(259*4)+3] <= 1'b0;
                  spc259_inst_done         <= 0;
                  spc259_phy_pc_w          <= 0;
                end else begin
                  active_thread[(259*4)]   <= 1'b1;
                  active_thread[(259*4)+1] <= 1'b1;
                  active_thread[(259*4)+2] <= 1'b1;
                  active_thread[(259*4)+3] <= 1'b1;
                  spc259_inst_done         <= `ARIANE_CORE259.piton_pc_vld;
                  spc259_phy_pc_w          <= `ARIANE_CORE259.piton_pc;
                end
            end
    

            assign spc260_thread_id = 2'b00;
            assign spc260_rtl_pc = spc260_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(260*4)]   <= 1'b0;
                  active_thread[(260*4)+1] <= 1'b0;
                  active_thread[(260*4)+2] <= 1'b0;
                  active_thread[(260*4)+3] <= 1'b0;
                  spc260_inst_done         <= 0;
                  spc260_phy_pc_w          <= 0;
                end else begin
                  active_thread[(260*4)]   <= 1'b1;
                  active_thread[(260*4)+1] <= 1'b1;
                  active_thread[(260*4)+2] <= 1'b1;
                  active_thread[(260*4)+3] <= 1'b1;
                  spc260_inst_done         <= `ARIANE_CORE260.piton_pc_vld;
                  spc260_phy_pc_w          <= `ARIANE_CORE260.piton_pc;
                end
            end
    

            assign spc261_thread_id = 2'b00;
            assign spc261_rtl_pc = spc261_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(261*4)]   <= 1'b0;
                  active_thread[(261*4)+1] <= 1'b0;
                  active_thread[(261*4)+2] <= 1'b0;
                  active_thread[(261*4)+3] <= 1'b0;
                  spc261_inst_done         <= 0;
                  spc261_phy_pc_w          <= 0;
                end else begin
                  active_thread[(261*4)]   <= 1'b1;
                  active_thread[(261*4)+1] <= 1'b1;
                  active_thread[(261*4)+2] <= 1'b1;
                  active_thread[(261*4)+3] <= 1'b1;
                  spc261_inst_done         <= `ARIANE_CORE261.piton_pc_vld;
                  spc261_phy_pc_w          <= `ARIANE_CORE261.piton_pc;
                end
            end
    

            assign spc262_thread_id = 2'b00;
            assign spc262_rtl_pc = spc262_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(262*4)]   <= 1'b0;
                  active_thread[(262*4)+1] <= 1'b0;
                  active_thread[(262*4)+2] <= 1'b0;
                  active_thread[(262*4)+3] <= 1'b0;
                  spc262_inst_done         <= 0;
                  spc262_phy_pc_w          <= 0;
                end else begin
                  active_thread[(262*4)]   <= 1'b1;
                  active_thread[(262*4)+1] <= 1'b1;
                  active_thread[(262*4)+2] <= 1'b1;
                  active_thread[(262*4)+3] <= 1'b1;
                  spc262_inst_done         <= `ARIANE_CORE262.piton_pc_vld;
                  spc262_phy_pc_w          <= `ARIANE_CORE262.piton_pc;
                end
            end
    

            assign spc263_thread_id = 2'b00;
            assign spc263_rtl_pc = spc263_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(263*4)]   <= 1'b0;
                  active_thread[(263*4)+1] <= 1'b0;
                  active_thread[(263*4)+2] <= 1'b0;
                  active_thread[(263*4)+3] <= 1'b0;
                  spc263_inst_done         <= 0;
                  spc263_phy_pc_w          <= 0;
                end else begin
                  active_thread[(263*4)]   <= 1'b1;
                  active_thread[(263*4)+1] <= 1'b1;
                  active_thread[(263*4)+2] <= 1'b1;
                  active_thread[(263*4)+3] <= 1'b1;
                  spc263_inst_done         <= `ARIANE_CORE263.piton_pc_vld;
                  spc263_phy_pc_w          <= `ARIANE_CORE263.piton_pc;
                end
            end
    

            assign spc264_thread_id = 2'b00;
            assign spc264_rtl_pc = spc264_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(264*4)]   <= 1'b0;
                  active_thread[(264*4)+1] <= 1'b0;
                  active_thread[(264*4)+2] <= 1'b0;
                  active_thread[(264*4)+3] <= 1'b0;
                  spc264_inst_done         <= 0;
                  spc264_phy_pc_w          <= 0;
                end else begin
                  active_thread[(264*4)]   <= 1'b1;
                  active_thread[(264*4)+1] <= 1'b1;
                  active_thread[(264*4)+2] <= 1'b1;
                  active_thread[(264*4)+3] <= 1'b1;
                  spc264_inst_done         <= `ARIANE_CORE264.piton_pc_vld;
                  spc264_phy_pc_w          <= `ARIANE_CORE264.piton_pc;
                end
            end
    

            assign spc265_thread_id = 2'b00;
            assign spc265_rtl_pc = spc265_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(265*4)]   <= 1'b0;
                  active_thread[(265*4)+1] <= 1'b0;
                  active_thread[(265*4)+2] <= 1'b0;
                  active_thread[(265*4)+3] <= 1'b0;
                  spc265_inst_done         <= 0;
                  spc265_phy_pc_w          <= 0;
                end else begin
                  active_thread[(265*4)]   <= 1'b1;
                  active_thread[(265*4)+1] <= 1'b1;
                  active_thread[(265*4)+2] <= 1'b1;
                  active_thread[(265*4)+3] <= 1'b1;
                  spc265_inst_done         <= `ARIANE_CORE265.piton_pc_vld;
                  spc265_phy_pc_w          <= `ARIANE_CORE265.piton_pc;
                end
            end
    

            assign spc266_thread_id = 2'b00;
            assign spc266_rtl_pc = spc266_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(266*4)]   <= 1'b0;
                  active_thread[(266*4)+1] <= 1'b0;
                  active_thread[(266*4)+2] <= 1'b0;
                  active_thread[(266*4)+3] <= 1'b0;
                  spc266_inst_done         <= 0;
                  spc266_phy_pc_w          <= 0;
                end else begin
                  active_thread[(266*4)]   <= 1'b1;
                  active_thread[(266*4)+1] <= 1'b1;
                  active_thread[(266*4)+2] <= 1'b1;
                  active_thread[(266*4)+3] <= 1'b1;
                  spc266_inst_done         <= `ARIANE_CORE266.piton_pc_vld;
                  spc266_phy_pc_w          <= `ARIANE_CORE266.piton_pc;
                end
            end
    

            assign spc267_thread_id = 2'b00;
            assign spc267_rtl_pc = spc267_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(267*4)]   <= 1'b0;
                  active_thread[(267*4)+1] <= 1'b0;
                  active_thread[(267*4)+2] <= 1'b0;
                  active_thread[(267*4)+3] <= 1'b0;
                  spc267_inst_done         <= 0;
                  spc267_phy_pc_w          <= 0;
                end else begin
                  active_thread[(267*4)]   <= 1'b1;
                  active_thread[(267*4)+1] <= 1'b1;
                  active_thread[(267*4)+2] <= 1'b1;
                  active_thread[(267*4)+3] <= 1'b1;
                  spc267_inst_done         <= `ARIANE_CORE267.piton_pc_vld;
                  spc267_phy_pc_w          <= `ARIANE_CORE267.piton_pc;
                end
            end
    

            assign spc268_thread_id = 2'b00;
            assign spc268_rtl_pc = spc268_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(268*4)]   <= 1'b0;
                  active_thread[(268*4)+1] <= 1'b0;
                  active_thread[(268*4)+2] <= 1'b0;
                  active_thread[(268*4)+3] <= 1'b0;
                  spc268_inst_done         <= 0;
                  spc268_phy_pc_w          <= 0;
                end else begin
                  active_thread[(268*4)]   <= 1'b1;
                  active_thread[(268*4)+1] <= 1'b1;
                  active_thread[(268*4)+2] <= 1'b1;
                  active_thread[(268*4)+3] <= 1'b1;
                  spc268_inst_done         <= `ARIANE_CORE268.piton_pc_vld;
                  spc268_phy_pc_w          <= `ARIANE_CORE268.piton_pc;
                end
            end
    

            assign spc269_thread_id = 2'b00;
            assign spc269_rtl_pc = spc269_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(269*4)]   <= 1'b0;
                  active_thread[(269*4)+1] <= 1'b0;
                  active_thread[(269*4)+2] <= 1'b0;
                  active_thread[(269*4)+3] <= 1'b0;
                  spc269_inst_done         <= 0;
                  spc269_phy_pc_w          <= 0;
                end else begin
                  active_thread[(269*4)]   <= 1'b1;
                  active_thread[(269*4)+1] <= 1'b1;
                  active_thread[(269*4)+2] <= 1'b1;
                  active_thread[(269*4)+3] <= 1'b1;
                  spc269_inst_done         <= `ARIANE_CORE269.piton_pc_vld;
                  spc269_phy_pc_w          <= `ARIANE_CORE269.piton_pc;
                end
            end
    

            assign spc270_thread_id = 2'b00;
            assign spc270_rtl_pc = spc270_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(270*4)]   <= 1'b0;
                  active_thread[(270*4)+1] <= 1'b0;
                  active_thread[(270*4)+2] <= 1'b0;
                  active_thread[(270*4)+3] <= 1'b0;
                  spc270_inst_done         <= 0;
                  spc270_phy_pc_w          <= 0;
                end else begin
                  active_thread[(270*4)]   <= 1'b1;
                  active_thread[(270*4)+1] <= 1'b1;
                  active_thread[(270*4)+2] <= 1'b1;
                  active_thread[(270*4)+3] <= 1'b1;
                  spc270_inst_done         <= `ARIANE_CORE270.piton_pc_vld;
                  spc270_phy_pc_w          <= `ARIANE_CORE270.piton_pc;
                end
            end
    

            assign spc271_thread_id = 2'b00;
            assign spc271_rtl_pc = spc271_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(271*4)]   <= 1'b0;
                  active_thread[(271*4)+1] <= 1'b0;
                  active_thread[(271*4)+2] <= 1'b0;
                  active_thread[(271*4)+3] <= 1'b0;
                  spc271_inst_done         <= 0;
                  spc271_phy_pc_w          <= 0;
                end else begin
                  active_thread[(271*4)]   <= 1'b1;
                  active_thread[(271*4)+1] <= 1'b1;
                  active_thread[(271*4)+2] <= 1'b1;
                  active_thread[(271*4)+3] <= 1'b1;
                  spc271_inst_done         <= `ARIANE_CORE271.piton_pc_vld;
                  spc271_phy_pc_w          <= `ARIANE_CORE271.piton_pc;
                end
            end
    

            assign spc272_thread_id = 2'b00;
            assign spc272_rtl_pc = spc272_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(272*4)]   <= 1'b0;
                  active_thread[(272*4)+1] <= 1'b0;
                  active_thread[(272*4)+2] <= 1'b0;
                  active_thread[(272*4)+3] <= 1'b0;
                  spc272_inst_done         <= 0;
                  spc272_phy_pc_w          <= 0;
                end else begin
                  active_thread[(272*4)]   <= 1'b1;
                  active_thread[(272*4)+1] <= 1'b1;
                  active_thread[(272*4)+2] <= 1'b1;
                  active_thread[(272*4)+3] <= 1'b1;
                  spc272_inst_done         <= `ARIANE_CORE272.piton_pc_vld;
                  spc272_phy_pc_w          <= `ARIANE_CORE272.piton_pc;
                end
            end
    

            assign spc273_thread_id = 2'b00;
            assign spc273_rtl_pc = spc273_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(273*4)]   <= 1'b0;
                  active_thread[(273*4)+1] <= 1'b0;
                  active_thread[(273*4)+2] <= 1'b0;
                  active_thread[(273*4)+3] <= 1'b0;
                  spc273_inst_done         <= 0;
                  spc273_phy_pc_w          <= 0;
                end else begin
                  active_thread[(273*4)]   <= 1'b1;
                  active_thread[(273*4)+1] <= 1'b1;
                  active_thread[(273*4)+2] <= 1'b1;
                  active_thread[(273*4)+3] <= 1'b1;
                  spc273_inst_done         <= `ARIANE_CORE273.piton_pc_vld;
                  spc273_phy_pc_w          <= `ARIANE_CORE273.piton_pc;
                end
            end
    

            assign spc274_thread_id = 2'b00;
            assign spc274_rtl_pc = spc274_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(274*4)]   <= 1'b0;
                  active_thread[(274*4)+1] <= 1'b0;
                  active_thread[(274*4)+2] <= 1'b0;
                  active_thread[(274*4)+3] <= 1'b0;
                  spc274_inst_done         <= 0;
                  spc274_phy_pc_w          <= 0;
                end else begin
                  active_thread[(274*4)]   <= 1'b1;
                  active_thread[(274*4)+1] <= 1'b1;
                  active_thread[(274*4)+2] <= 1'b1;
                  active_thread[(274*4)+3] <= 1'b1;
                  spc274_inst_done         <= `ARIANE_CORE274.piton_pc_vld;
                  spc274_phy_pc_w          <= `ARIANE_CORE274.piton_pc;
                end
            end
    

            assign spc275_thread_id = 2'b00;
            assign spc275_rtl_pc = spc275_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(275*4)]   <= 1'b0;
                  active_thread[(275*4)+1] <= 1'b0;
                  active_thread[(275*4)+2] <= 1'b0;
                  active_thread[(275*4)+3] <= 1'b0;
                  spc275_inst_done         <= 0;
                  spc275_phy_pc_w          <= 0;
                end else begin
                  active_thread[(275*4)]   <= 1'b1;
                  active_thread[(275*4)+1] <= 1'b1;
                  active_thread[(275*4)+2] <= 1'b1;
                  active_thread[(275*4)+3] <= 1'b1;
                  spc275_inst_done         <= `ARIANE_CORE275.piton_pc_vld;
                  spc275_phy_pc_w          <= `ARIANE_CORE275.piton_pc;
                end
            end
    

            assign spc276_thread_id = 2'b00;
            assign spc276_rtl_pc = spc276_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(276*4)]   <= 1'b0;
                  active_thread[(276*4)+1] <= 1'b0;
                  active_thread[(276*4)+2] <= 1'b0;
                  active_thread[(276*4)+3] <= 1'b0;
                  spc276_inst_done         <= 0;
                  spc276_phy_pc_w          <= 0;
                end else begin
                  active_thread[(276*4)]   <= 1'b1;
                  active_thread[(276*4)+1] <= 1'b1;
                  active_thread[(276*4)+2] <= 1'b1;
                  active_thread[(276*4)+3] <= 1'b1;
                  spc276_inst_done         <= `ARIANE_CORE276.piton_pc_vld;
                  spc276_phy_pc_w          <= `ARIANE_CORE276.piton_pc;
                end
            end
    

            assign spc277_thread_id = 2'b00;
            assign spc277_rtl_pc = spc277_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(277*4)]   <= 1'b0;
                  active_thread[(277*4)+1] <= 1'b0;
                  active_thread[(277*4)+2] <= 1'b0;
                  active_thread[(277*4)+3] <= 1'b0;
                  spc277_inst_done         <= 0;
                  spc277_phy_pc_w          <= 0;
                end else begin
                  active_thread[(277*4)]   <= 1'b1;
                  active_thread[(277*4)+1] <= 1'b1;
                  active_thread[(277*4)+2] <= 1'b1;
                  active_thread[(277*4)+3] <= 1'b1;
                  spc277_inst_done         <= `ARIANE_CORE277.piton_pc_vld;
                  spc277_phy_pc_w          <= `ARIANE_CORE277.piton_pc;
                end
            end
    

            assign spc278_thread_id = 2'b00;
            assign spc278_rtl_pc = spc278_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(278*4)]   <= 1'b0;
                  active_thread[(278*4)+1] <= 1'b0;
                  active_thread[(278*4)+2] <= 1'b0;
                  active_thread[(278*4)+3] <= 1'b0;
                  spc278_inst_done         <= 0;
                  spc278_phy_pc_w          <= 0;
                end else begin
                  active_thread[(278*4)]   <= 1'b1;
                  active_thread[(278*4)+1] <= 1'b1;
                  active_thread[(278*4)+2] <= 1'b1;
                  active_thread[(278*4)+3] <= 1'b1;
                  spc278_inst_done         <= `ARIANE_CORE278.piton_pc_vld;
                  spc278_phy_pc_w          <= `ARIANE_CORE278.piton_pc;
                end
            end
    

            assign spc279_thread_id = 2'b00;
            assign spc279_rtl_pc = spc279_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(279*4)]   <= 1'b0;
                  active_thread[(279*4)+1] <= 1'b0;
                  active_thread[(279*4)+2] <= 1'b0;
                  active_thread[(279*4)+3] <= 1'b0;
                  spc279_inst_done         <= 0;
                  spc279_phy_pc_w          <= 0;
                end else begin
                  active_thread[(279*4)]   <= 1'b1;
                  active_thread[(279*4)+1] <= 1'b1;
                  active_thread[(279*4)+2] <= 1'b1;
                  active_thread[(279*4)+3] <= 1'b1;
                  spc279_inst_done         <= `ARIANE_CORE279.piton_pc_vld;
                  spc279_phy_pc_w          <= `ARIANE_CORE279.piton_pc;
                end
            end
    

            assign spc280_thread_id = 2'b00;
            assign spc280_rtl_pc = spc280_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(280*4)]   <= 1'b0;
                  active_thread[(280*4)+1] <= 1'b0;
                  active_thread[(280*4)+2] <= 1'b0;
                  active_thread[(280*4)+3] <= 1'b0;
                  spc280_inst_done         <= 0;
                  spc280_phy_pc_w          <= 0;
                end else begin
                  active_thread[(280*4)]   <= 1'b1;
                  active_thread[(280*4)+1] <= 1'b1;
                  active_thread[(280*4)+2] <= 1'b1;
                  active_thread[(280*4)+3] <= 1'b1;
                  spc280_inst_done         <= `ARIANE_CORE280.piton_pc_vld;
                  spc280_phy_pc_w          <= `ARIANE_CORE280.piton_pc;
                end
            end
    

            assign spc281_thread_id = 2'b00;
            assign spc281_rtl_pc = spc281_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(281*4)]   <= 1'b0;
                  active_thread[(281*4)+1] <= 1'b0;
                  active_thread[(281*4)+2] <= 1'b0;
                  active_thread[(281*4)+3] <= 1'b0;
                  spc281_inst_done         <= 0;
                  spc281_phy_pc_w          <= 0;
                end else begin
                  active_thread[(281*4)]   <= 1'b1;
                  active_thread[(281*4)+1] <= 1'b1;
                  active_thread[(281*4)+2] <= 1'b1;
                  active_thread[(281*4)+3] <= 1'b1;
                  spc281_inst_done         <= `ARIANE_CORE281.piton_pc_vld;
                  spc281_phy_pc_w          <= `ARIANE_CORE281.piton_pc;
                end
            end
    

            assign spc282_thread_id = 2'b00;
            assign spc282_rtl_pc = spc282_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(282*4)]   <= 1'b0;
                  active_thread[(282*4)+1] <= 1'b0;
                  active_thread[(282*4)+2] <= 1'b0;
                  active_thread[(282*4)+3] <= 1'b0;
                  spc282_inst_done         <= 0;
                  spc282_phy_pc_w          <= 0;
                end else begin
                  active_thread[(282*4)]   <= 1'b1;
                  active_thread[(282*4)+1] <= 1'b1;
                  active_thread[(282*4)+2] <= 1'b1;
                  active_thread[(282*4)+3] <= 1'b1;
                  spc282_inst_done         <= `ARIANE_CORE282.piton_pc_vld;
                  spc282_phy_pc_w          <= `ARIANE_CORE282.piton_pc;
                end
            end
    

            assign spc283_thread_id = 2'b00;
            assign spc283_rtl_pc = spc283_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(283*4)]   <= 1'b0;
                  active_thread[(283*4)+1] <= 1'b0;
                  active_thread[(283*4)+2] <= 1'b0;
                  active_thread[(283*4)+3] <= 1'b0;
                  spc283_inst_done         <= 0;
                  spc283_phy_pc_w          <= 0;
                end else begin
                  active_thread[(283*4)]   <= 1'b1;
                  active_thread[(283*4)+1] <= 1'b1;
                  active_thread[(283*4)+2] <= 1'b1;
                  active_thread[(283*4)+3] <= 1'b1;
                  spc283_inst_done         <= `ARIANE_CORE283.piton_pc_vld;
                  spc283_phy_pc_w          <= `ARIANE_CORE283.piton_pc;
                end
            end
    

            assign spc284_thread_id = 2'b00;
            assign spc284_rtl_pc = spc284_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(284*4)]   <= 1'b0;
                  active_thread[(284*4)+1] <= 1'b0;
                  active_thread[(284*4)+2] <= 1'b0;
                  active_thread[(284*4)+3] <= 1'b0;
                  spc284_inst_done         <= 0;
                  spc284_phy_pc_w          <= 0;
                end else begin
                  active_thread[(284*4)]   <= 1'b1;
                  active_thread[(284*4)+1] <= 1'b1;
                  active_thread[(284*4)+2] <= 1'b1;
                  active_thread[(284*4)+3] <= 1'b1;
                  spc284_inst_done         <= `ARIANE_CORE284.piton_pc_vld;
                  spc284_phy_pc_w          <= `ARIANE_CORE284.piton_pc;
                end
            end
    

            assign spc285_thread_id = 2'b00;
            assign spc285_rtl_pc = spc285_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(285*4)]   <= 1'b0;
                  active_thread[(285*4)+1] <= 1'b0;
                  active_thread[(285*4)+2] <= 1'b0;
                  active_thread[(285*4)+3] <= 1'b0;
                  spc285_inst_done         <= 0;
                  spc285_phy_pc_w          <= 0;
                end else begin
                  active_thread[(285*4)]   <= 1'b1;
                  active_thread[(285*4)+1] <= 1'b1;
                  active_thread[(285*4)+2] <= 1'b1;
                  active_thread[(285*4)+3] <= 1'b1;
                  spc285_inst_done         <= `ARIANE_CORE285.piton_pc_vld;
                  spc285_phy_pc_w          <= `ARIANE_CORE285.piton_pc;
                end
            end
    

            assign spc286_thread_id = 2'b00;
            assign spc286_rtl_pc = spc286_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(286*4)]   <= 1'b0;
                  active_thread[(286*4)+1] <= 1'b0;
                  active_thread[(286*4)+2] <= 1'b0;
                  active_thread[(286*4)+3] <= 1'b0;
                  spc286_inst_done         <= 0;
                  spc286_phy_pc_w          <= 0;
                end else begin
                  active_thread[(286*4)]   <= 1'b1;
                  active_thread[(286*4)+1] <= 1'b1;
                  active_thread[(286*4)+2] <= 1'b1;
                  active_thread[(286*4)+3] <= 1'b1;
                  spc286_inst_done         <= `ARIANE_CORE286.piton_pc_vld;
                  spc286_phy_pc_w          <= `ARIANE_CORE286.piton_pc;
                end
            end
    

            assign spc287_thread_id = 2'b00;
            assign spc287_rtl_pc = spc287_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(287*4)]   <= 1'b0;
                  active_thread[(287*4)+1] <= 1'b0;
                  active_thread[(287*4)+2] <= 1'b0;
                  active_thread[(287*4)+3] <= 1'b0;
                  spc287_inst_done         <= 0;
                  spc287_phy_pc_w          <= 0;
                end else begin
                  active_thread[(287*4)]   <= 1'b1;
                  active_thread[(287*4)+1] <= 1'b1;
                  active_thread[(287*4)+2] <= 1'b1;
                  active_thread[(287*4)+3] <= 1'b1;
                  spc287_inst_done         <= `ARIANE_CORE287.piton_pc_vld;
                  spc287_phy_pc_w          <= `ARIANE_CORE287.piton_pc;
                end
            end
    

            assign spc288_thread_id = 2'b00;
            assign spc288_rtl_pc = spc288_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(288*4)]   <= 1'b0;
                  active_thread[(288*4)+1] <= 1'b0;
                  active_thread[(288*4)+2] <= 1'b0;
                  active_thread[(288*4)+3] <= 1'b0;
                  spc288_inst_done         <= 0;
                  spc288_phy_pc_w          <= 0;
                end else begin
                  active_thread[(288*4)]   <= 1'b1;
                  active_thread[(288*4)+1] <= 1'b1;
                  active_thread[(288*4)+2] <= 1'b1;
                  active_thread[(288*4)+3] <= 1'b1;
                  spc288_inst_done         <= `ARIANE_CORE288.piton_pc_vld;
                  spc288_phy_pc_w          <= `ARIANE_CORE288.piton_pc;
                end
            end
    

            assign spc289_thread_id = 2'b00;
            assign spc289_rtl_pc = spc289_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(289*4)]   <= 1'b0;
                  active_thread[(289*4)+1] <= 1'b0;
                  active_thread[(289*4)+2] <= 1'b0;
                  active_thread[(289*4)+3] <= 1'b0;
                  spc289_inst_done         <= 0;
                  spc289_phy_pc_w          <= 0;
                end else begin
                  active_thread[(289*4)]   <= 1'b1;
                  active_thread[(289*4)+1] <= 1'b1;
                  active_thread[(289*4)+2] <= 1'b1;
                  active_thread[(289*4)+3] <= 1'b1;
                  spc289_inst_done         <= `ARIANE_CORE289.piton_pc_vld;
                  spc289_phy_pc_w          <= `ARIANE_CORE289.piton_pc;
                end
            end
    

            assign spc290_thread_id = 2'b00;
            assign spc290_rtl_pc = spc290_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(290*4)]   <= 1'b0;
                  active_thread[(290*4)+1] <= 1'b0;
                  active_thread[(290*4)+2] <= 1'b0;
                  active_thread[(290*4)+3] <= 1'b0;
                  spc290_inst_done         <= 0;
                  spc290_phy_pc_w          <= 0;
                end else begin
                  active_thread[(290*4)]   <= 1'b1;
                  active_thread[(290*4)+1] <= 1'b1;
                  active_thread[(290*4)+2] <= 1'b1;
                  active_thread[(290*4)+3] <= 1'b1;
                  spc290_inst_done         <= `ARIANE_CORE290.piton_pc_vld;
                  spc290_phy_pc_w          <= `ARIANE_CORE290.piton_pc;
                end
            end
    

            assign spc291_thread_id = 2'b00;
            assign spc291_rtl_pc = spc291_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(291*4)]   <= 1'b0;
                  active_thread[(291*4)+1] <= 1'b0;
                  active_thread[(291*4)+2] <= 1'b0;
                  active_thread[(291*4)+3] <= 1'b0;
                  spc291_inst_done         <= 0;
                  spc291_phy_pc_w          <= 0;
                end else begin
                  active_thread[(291*4)]   <= 1'b1;
                  active_thread[(291*4)+1] <= 1'b1;
                  active_thread[(291*4)+2] <= 1'b1;
                  active_thread[(291*4)+3] <= 1'b1;
                  spc291_inst_done         <= `ARIANE_CORE291.piton_pc_vld;
                  spc291_phy_pc_w          <= `ARIANE_CORE291.piton_pc;
                end
            end
    

            assign spc292_thread_id = 2'b00;
            assign spc292_rtl_pc = spc292_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(292*4)]   <= 1'b0;
                  active_thread[(292*4)+1] <= 1'b0;
                  active_thread[(292*4)+2] <= 1'b0;
                  active_thread[(292*4)+3] <= 1'b0;
                  spc292_inst_done         <= 0;
                  spc292_phy_pc_w          <= 0;
                end else begin
                  active_thread[(292*4)]   <= 1'b1;
                  active_thread[(292*4)+1] <= 1'b1;
                  active_thread[(292*4)+2] <= 1'b1;
                  active_thread[(292*4)+3] <= 1'b1;
                  spc292_inst_done         <= `ARIANE_CORE292.piton_pc_vld;
                  spc292_phy_pc_w          <= `ARIANE_CORE292.piton_pc;
                end
            end
    

            assign spc293_thread_id = 2'b00;
            assign spc293_rtl_pc = spc293_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(293*4)]   <= 1'b0;
                  active_thread[(293*4)+1] <= 1'b0;
                  active_thread[(293*4)+2] <= 1'b0;
                  active_thread[(293*4)+3] <= 1'b0;
                  spc293_inst_done         <= 0;
                  spc293_phy_pc_w          <= 0;
                end else begin
                  active_thread[(293*4)]   <= 1'b1;
                  active_thread[(293*4)+1] <= 1'b1;
                  active_thread[(293*4)+2] <= 1'b1;
                  active_thread[(293*4)+3] <= 1'b1;
                  spc293_inst_done         <= `ARIANE_CORE293.piton_pc_vld;
                  spc293_phy_pc_w          <= `ARIANE_CORE293.piton_pc;
                end
            end
    

            assign spc294_thread_id = 2'b00;
            assign spc294_rtl_pc = spc294_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(294*4)]   <= 1'b0;
                  active_thread[(294*4)+1] <= 1'b0;
                  active_thread[(294*4)+2] <= 1'b0;
                  active_thread[(294*4)+3] <= 1'b0;
                  spc294_inst_done         <= 0;
                  spc294_phy_pc_w          <= 0;
                end else begin
                  active_thread[(294*4)]   <= 1'b1;
                  active_thread[(294*4)+1] <= 1'b1;
                  active_thread[(294*4)+2] <= 1'b1;
                  active_thread[(294*4)+3] <= 1'b1;
                  spc294_inst_done         <= `ARIANE_CORE294.piton_pc_vld;
                  spc294_phy_pc_w          <= `ARIANE_CORE294.piton_pc;
                end
            end
    

            assign spc295_thread_id = 2'b00;
            assign spc295_rtl_pc = spc295_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(295*4)]   <= 1'b0;
                  active_thread[(295*4)+1] <= 1'b0;
                  active_thread[(295*4)+2] <= 1'b0;
                  active_thread[(295*4)+3] <= 1'b0;
                  spc295_inst_done         <= 0;
                  spc295_phy_pc_w          <= 0;
                end else begin
                  active_thread[(295*4)]   <= 1'b1;
                  active_thread[(295*4)+1] <= 1'b1;
                  active_thread[(295*4)+2] <= 1'b1;
                  active_thread[(295*4)+3] <= 1'b1;
                  spc295_inst_done         <= `ARIANE_CORE295.piton_pc_vld;
                  spc295_phy_pc_w          <= `ARIANE_CORE295.piton_pc;
                end
            end
    

            assign spc296_thread_id = 2'b00;
            assign spc296_rtl_pc = spc296_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(296*4)]   <= 1'b0;
                  active_thread[(296*4)+1] <= 1'b0;
                  active_thread[(296*4)+2] <= 1'b0;
                  active_thread[(296*4)+3] <= 1'b0;
                  spc296_inst_done         <= 0;
                  spc296_phy_pc_w          <= 0;
                end else begin
                  active_thread[(296*4)]   <= 1'b1;
                  active_thread[(296*4)+1] <= 1'b1;
                  active_thread[(296*4)+2] <= 1'b1;
                  active_thread[(296*4)+3] <= 1'b1;
                  spc296_inst_done         <= `ARIANE_CORE296.piton_pc_vld;
                  spc296_phy_pc_w          <= `ARIANE_CORE296.piton_pc;
                end
            end
    

            assign spc297_thread_id = 2'b00;
            assign spc297_rtl_pc = spc297_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(297*4)]   <= 1'b0;
                  active_thread[(297*4)+1] <= 1'b0;
                  active_thread[(297*4)+2] <= 1'b0;
                  active_thread[(297*4)+3] <= 1'b0;
                  spc297_inst_done         <= 0;
                  spc297_phy_pc_w          <= 0;
                end else begin
                  active_thread[(297*4)]   <= 1'b1;
                  active_thread[(297*4)+1] <= 1'b1;
                  active_thread[(297*4)+2] <= 1'b1;
                  active_thread[(297*4)+3] <= 1'b1;
                  spc297_inst_done         <= `ARIANE_CORE297.piton_pc_vld;
                  spc297_phy_pc_w          <= `ARIANE_CORE297.piton_pc;
                end
            end
    

            assign spc298_thread_id = 2'b00;
            assign spc298_rtl_pc = spc298_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(298*4)]   <= 1'b0;
                  active_thread[(298*4)+1] <= 1'b0;
                  active_thread[(298*4)+2] <= 1'b0;
                  active_thread[(298*4)+3] <= 1'b0;
                  spc298_inst_done         <= 0;
                  spc298_phy_pc_w          <= 0;
                end else begin
                  active_thread[(298*4)]   <= 1'b1;
                  active_thread[(298*4)+1] <= 1'b1;
                  active_thread[(298*4)+2] <= 1'b1;
                  active_thread[(298*4)+3] <= 1'b1;
                  spc298_inst_done         <= `ARIANE_CORE298.piton_pc_vld;
                  spc298_phy_pc_w          <= `ARIANE_CORE298.piton_pc;
                end
            end
    

            assign spc299_thread_id = 2'b00;
            assign spc299_rtl_pc = spc299_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(299*4)]   <= 1'b0;
                  active_thread[(299*4)+1] <= 1'b0;
                  active_thread[(299*4)+2] <= 1'b0;
                  active_thread[(299*4)+3] <= 1'b0;
                  spc299_inst_done         <= 0;
                  spc299_phy_pc_w          <= 0;
                end else begin
                  active_thread[(299*4)]   <= 1'b1;
                  active_thread[(299*4)+1] <= 1'b1;
                  active_thread[(299*4)+2] <= 1'b1;
                  active_thread[(299*4)+3] <= 1'b1;
                  spc299_inst_done         <= `ARIANE_CORE299.piton_pc_vld;
                  spc299_phy_pc_w          <= `ARIANE_CORE299.piton_pc;
                end
            end
    

            assign spc300_thread_id = 2'b00;
            assign spc300_rtl_pc = spc300_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(300*4)]   <= 1'b0;
                  active_thread[(300*4)+1] <= 1'b0;
                  active_thread[(300*4)+2] <= 1'b0;
                  active_thread[(300*4)+3] <= 1'b0;
                  spc300_inst_done         <= 0;
                  spc300_phy_pc_w          <= 0;
                end else begin
                  active_thread[(300*4)]   <= 1'b1;
                  active_thread[(300*4)+1] <= 1'b1;
                  active_thread[(300*4)+2] <= 1'b1;
                  active_thread[(300*4)+3] <= 1'b1;
                  spc300_inst_done         <= `ARIANE_CORE300.piton_pc_vld;
                  spc300_phy_pc_w          <= `ARIANE_CORE300.piton_pc;
                end
            end
    

            assign spc301_thread_id = 2'b00;
            assign spc301_rtl_pc = spc301_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(301*4)]   <= 1'b0;
                  active_thread[(301*4)+1] <= 1'b0;
                  active_thread[(301*4)+2] <= 1'b0;
                  active_thread[(301*4)+3] <= 1'b0;
                  spc301_inst_done         <= 0;
                  spc301_phy_pc_w          <= 0;
                end else begin
                  active_thread[(301*4)]   <= 1'b1;
                  active_thread[(301*4)+1] <= 1'b1;
                  active_thread[(301*4)+2] <= 1'b1;
                  active_thread[(301*4)+3] <= 1'b1;
                  spc301_inst_done         <= `ARIANE_CORE301.piton_pc_vld;
                  spc301_phy_pc_w          <= `ARIANE_CORE301.piton_pc;
                end
            end
    

            assign spc302_thread_id = 2'b00;
            assign spc302_rtl_pc = spc302_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(302*4)]   <= 1'b0;
                  active_thread[(302*4)+1] <= 1'b0;
                  active_thread[(302*4)+2] <= 1'b0;
                  active_thread[(302*4)+3] <= 1'b0;
                  spc302_inst_done         <= 0;
                  spc302_phy_pc_w          <= 0;
                end else begin
                  active_thread[(302*4)]   <= 1'b1;
                  active_thread[(302*4)+1] <= 1'b1;
                  active_thread[(302*4)+2] <= 1'b1;
                  active_thread[(302*4)+3] <= 1'b1;
                  spc302_inst_done         <= `ARIANE_CORE302.piton_pc_vld;
                  spc302_phy_pc_w          <= `ARIANE_CORE302.piton_pc;
                end
            end
    

            assign spc303_thread_id = 2'b00;
            assign spc303_rtl_pc = spc303_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(303*4)]   <= 1'b0;
                  active_thread[(303*4)+1] <= 1'b0;
                  active_thread[(303*4)+2] <= 1'b0;
                  active_thread[(303*4)+3] <= 1'b0;
                  spc303_inst_done         <= 0;
                  spc303_phy_pc_w          <= 0;
                end else begin
                  active_thread[(303*4)]   <= 1'b1;
                  active_thread[(303*4)+1] <= 1'b1;
                  active_thread[(303*4)+2] <= 1'b1;
                  active_thread[(303*4)+3] <= 1'b1;
                  spc303_inst_done         <= `ARIANE_CORE303.piton_pc_vld;
                  spc303_phy_pc_w          <= `ARIANE_CORE303.piton_pc;
                end
            end
    

            assign spc304_thread_id = 2'b00;
            assign spc304_rtl_pc = spc304_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(304*4)]   <= 1'b0;
                  active_thread[(304*4)+1] <= 1'b0;
                  active_thread[(304*4)+2] <= 1'b0;
                  active_thread[(304*4)+3] <= 1'b0;
                  spc304_inst_done         <= 0;
                  spc304_phy_pc_w          <= 0;
                end else begin
                  active_thread[(304*4)]   <= 1'b1;
                  active_thread[(304*4)+1] <= 1'b1;
                  active_thread[(304*4)+2] <= 1'b1;
                  active_thread[(304*4)+3] <= 1'b1;
                  spc304_inst_done         <= `ARIANE_CORE304.piton_pc_vld;
                  spc304_phy_pc_w          <= `ARIANE_CORE304.piton_pc;
                end
            end
    

            assign spc305_thread_id = 2'b00;
            assign spc305_rtl_pc = spc305_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(305*4)]   <= 1'b0;
                  active_thread[(305*4)+1] <= 1'b0;
                  active_thread[(305*4)+2] <= 1'b0;
                  active_thread[(305*4)+3] <= 1'b0;
                  spc305_inst_done         <= 0;
                  spc305_phy_pc_w          <= 0;
                end else begin
                  active_thread[(305*4)]   <= 1'b1;
                  active_thread[(305*4)+1] <= 1'b1;
                  active_thread[(305*4)+2] <= 1'b1;
                  active_thread[(305*4)+3] <= 1'b1;
                  spc305_inst_done         <= `ARIANE_CORE305.piton_pc_vld;
                  spc305_phy_pc_w          <= `ARIANE_CORE305.piton_pc;
                end
            end
    

            assign spc306_thread_id = 2'b00;
            assign spc306_rtl_pc = spc306_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(306*4)]   <= 1'b0;
                  active_thread[(306*4)+1] <= 1'b0;
                  active_thread[(306*4)+2] <= 1'b0;
                  active_thread[(306*4)+3] <= 1'b0;
                  spc306_inst_done         <= 0;
                  spc306_phy_pc_w          <= 0;
                end else begin
                  active_thread[(306*4)]   <= 1'b1;
                  active_thread[(306*4)+1] <= 1'b1;
                  active_thread[(306*4)+2] <= 1'b1;
                  active_thread[(306*4)+3] <= 1'b1;
                  spc306_inst_done         <= `ARIANE_CORE306.piton_pc_vld;
                  spc306_phy_pc_w          <= `ARIANE_CORE306.piton_pc;
                end
            end
    

            assign spc307_thread_id = 2'b00;
            assign spc307_rtl_pc = spc307_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(307*4)]   <= 1'b0;
                  active_thread[(307*4)+1] <= 1'b0;
                  active_thread[(307*4)+2] <= 1'b0;
                  active_thread[(307*4)+3] <= 1'b0;
                  spc307_inst_done         <= 0;
                  spc307_phy_pc_w          <= 0;
                end else begin
                  active_thread[(307*4)]   <= 1'b1;
                  active_thread[(307*4)+1] <= 1'b1;
                  active_thread[(307*4)+2] <= 1'b1;
                  active_thread[(307*4)+3] <= 1'b1;
                  spc307_inst_done         <= `ARIANE_CORE307.piton_pc_vld;
                  spc307_phy_pc_w          <= `ARIANE_CORE307.piton_pc;
                end
            end
    

            assign spc308_thread_id = 2'b00;
            assign spc308_rtl_pc = spc308_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(308*4)]   <= 1'b0;
                  active_thread[(308*4)+1] <= 1'b0;
                  active_thread[(308*4)+2] <= 1'b0;
                  active_thread[(308*4)+3] <= 1'b0;
                  spc308_inst_done         <= 0;
                  spc308_phy_pc_w          <= 0;
                end else begin
                  active_thread[(308*4)]   <= 1'b1;
                  active_thread[(308*4)+1] <= 1'b1;
                  active_thread[(308*4)+2] <= 1'b1;
                  active_thread[(308*4)+3] <= 1'b1;
                  spc308_inst_done         <= `ARIANE_CORE308.piton_pc_vld;
                  spc308_phy_pc_w          <= `ARIANE_CORE308.piton_pc;
                end
            end
    

            assign spc309_thread_id = 2'b00;
            assign spc309_rtl_pc = spc309_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(309*4)]   <= 1'b0;
                  active_thread[(309*4)+1] <= 1'b0;
                  active_thread[(309*4)+2] <= 1'b0;
                  active_thread[(309*4)+3] <= 1'b0;
                  spc309_inst_done         <= 0;
                  spc309_phy_pc_w          <= 0;
                end else begin
                  active_thread[(309*4)]   <= 1'b1;
                  active_thread[(309*4)+1] <= 1'b1;
                  active_thread[(309*4)+2] <= 1'b1;
                  active_thread[(309*4)+3] <= 1'b1;
                  spc309_inst_done         <= `ARIANE_CORE309.piton_pc_vld;
                  spc309_phy_pc_w          <= `ARIANE_CORE309.piton_pc;
                end
            end
    

            assign spc310_thread_id = 2'b00;
            assign spc310_rtl_pc = spc310_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(310*4)]   <= 1'b0;
                  active_thread[(310*4)+1] <= 1'b0;
                  active_thread[(310*4)+2] <= 1'b0;
                  active_thread[(310*4)+3] <= 1'b0;
                  spc310_inst_done         <= 0;
                  spc310_phy_pc_w          <= 0;
                end else begin
                  active_thread[(310*4)]   <= 1'b1;
                  active_thread[(310*4)+1] <= 1'b1;
                  active_thread[(310*4)+2] <= 1'b1;
                  active_thread[(310*4)+3] <= 1'b1;
                  spc310_inst_done         <= `ARIANE_CORE310.piton_pc_vld;
                  spc310_phy_pc_w          <= `ARIANE_CORE310.piton_pc;
                end
            end
    

            assign spc311_thread_id = 2'b00;
            assign spc311_rtl_pc = spc311_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(311*4)]   <= 1'b0;
                  active_thread[(311*4)+1] <= 1'b0;
                  active_thread[(311*4)+2] <= 1'b0;
                  active_thread[(311*4)+3] <= 1'b0;
                  spc311_inst_done         <= 0;
                  spc311_phy_pc_w          <= 0;
                end else begin
                  active_thread[(311*4)]   <= 1'b1;
                  active_thread[(311*4)+1] <= 1'b1;
                  active_thread[(311*4)+2] <= 1'b1;
                  active_thread[(311*4)+3] <= 1'b1;
                  spc311_inst_done         <= `ARIANE_CORE311.piton_pc_vld;
                  spc311_phy_pc_w          <= `ARIANE_CORE311.piton_pc;
                end
            end
    

            assign spc312_thread_id = 2'b00;
            assign spc312_rtl_pc = spc312_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(312*4)]   <= 1'b0;
                  active_thread[(312*4)+1] <= 1'b0;
                  active_thread[(312*4)+2] <= 1'b0;
                  active_thread[(312*4)+3] <= 1'b0;
                  spc312_inst_done         <= 0;
                  spc312_phy_pc_w          <= 0;
                end else begin
                  active_thread[(312*4)]   <= 1'b1;
                  active_thread[(312*4)+1] <= 1'b1;
                  active_thread[(312*4)+2] <= 1'b1;
                  active_thread[(312*4)+3] <= 1'b1;
                  spc312_inst_done         <= `ARIANE_CORE312.piton_pc_vld;
                  spc312_phy_pc_w          <= `ARIANE_CORE312.piton_pc;
                end
            end
    

            assign spc313_thread_id = 2'b00;
            assign spc313_rtl_pc = spc313_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(313*4)]   <= 1'b0;
                  active_thread[(313*4)+1] <= 1'b0;
                  active_thread[(313*4)+2] <= 1'b0;
                  active_thread[(313*4)+3] <= 1'b0;
                  spc313_inst_done         <= 0;
                  spc313_phy_pc_w          <= 0;
                end else begin
                  active_thread[(313*4)]   <= 1'b1;
                  active_thread[(313*4)+1] <= 1'b1;
                  active_thread[(313*4)+2] <= 1'b1;
                  active_thread[(313*4)+3] <= 1'b1;
                  spc313_inst_done         <= `ARIANE_CORE313.piton_pc_vld;
                  spc313_phy_pc_w          <= `ARIANE_CORE313.piton_pc;
                end
            end
    

            assign spc314_thread_id = 2'b00;
            assign spc314_rtl_pc = spc314_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(314*4)]   <= 1'b0;
                  active_thread[(314*4)+1] <= 1'b0;
                  active_thread[(314*4)+2] <= 1'b0;
                  active_thread[(314*4)+3] <= 1'b0;
                  spc314_inst_done         <= 0;
                  spc314_phy_pc_w          <= 0;
                end else begin
                  active_thread[(314*4)]   <= 1'b1;
                  active_thread[(314*4)+1] <= 1'b1;
                  active_thread[(314*4)+2] <= 1'b1;
                  active_thread[(314*4)+3] <= 1'b1;
                  spc314_inst_done         <= `ARIANE_CORE314.piton_pc_vld;
                  spc314_phy_pc_w          <= `ARIANE_CORE314.piton_pc;
                end
            end
    

            assign spc315_thread_id = 2'b00;
            assign spc315_rtl_pc = spc315_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(315*4)]   <= 1'b0;
                  active_thread[(315*4)+1] <= 1'b0;
                  active_thread[(315*4)+2] <= 1'b0;
                  active_thread[(315*4)+3] <= 1'b0;
                  spc315_inst_done         <= 0;
                  spc315_phy_pc_w          <= 0;
                end else begin
                  active_thread[(315*4)]   <= 1'b1;
                  active_thread[(315*4)+1] <= 1'b1;
                  active_thread[(315*4)+2] <= 1'b1;
                  active_thread[(315*4)+3] <= 1'b1;
                  spc315_inst_done         <= `ARIANE_CORE315.piton_pc_vld;
                  spc315_phy_pc_w          <= `ARIANE_CORE315.piton_pc;
                end
            end
    

            assign spc316_thread_id = 2'b00;
            assign spc316_rtl_pc = spc316_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(316*4)]   <= 1'b0;
                  active_thread[(316*4)+1] <= 1'b0;
                  active_thread[(316*4)+2] <= 1'b0;
                  active_thread[(316*4)+3] <= 1'b0;
                  spc316_inst_done         <= 0;
                  spc316_phy_pc_w          <= 0;
                end else begin
                  active_thread[(316*4)]   <= 1'b1;
                  active_thread[(316*4)+1] <= 1'b1;
                  active_thread[(316*4)+2] <= 1'b1;
                  active_thread[(316*4)+3] <= 1'b1;
                  spc316_inst_done         <= `ARIANE_CORE316.piton_pc_vld;
                  spc316_phy_pc_w          <= `ARIANE_CORE316.piton_pc;
                end
            end
    

            assign spc317_thread_id = 2'b00;
            assign spc317_rtl_pc = spc317_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(317*4)]   <= 1'b0;
                  active_thread[(317*4)+1] <= 1'b0;
                  active_thread[(317*4)+2] <= 1'b0;
                  active_thread[(317*4)+3] <= 1'b0;
                  spc317_inst_done         <= 0;
                  spc317_phy_pc_w          <= 0;
                end else begin
                  active_thread[(317*4)]   <= 1'b1;
                  active_thread[(317*4)+1] <= 1'b1;
                  active_thread[(317*4)+2] <= 1'b1;
                  active_thread[(317*4)+3] <= 1'b1;
                  spc317_inst_done         <= `ARIANE_CORE317.piton_pc_vld;
                  spc317_phy_pc_w          <= `ARIANE_CORE317.piton_pc;
                end
            end
    

            assign spc318_thread_id = 2'b00;
            assign spc318_rtl_pc = spc318_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(318*4)]   <= 1'b0;
                  active_thread[(318*4)+1] <= 1'b0;
                  active_thread[(318*4)+2] <= 1'b0;
                  active_thread[(318*4)+3] <= 1'b0;
                  spc318_inst_done         <= 0;
                  spc318_phy_pc_w          <= 0;
                end else begin
                  active_thread[(318*4)]   <= 1'b1;
                  active_thread[(318*4)+1] <= 1'b1;
                  active_thread[(318*4)+2] <= 1'b1;
                  active_thread[(318*4)+3] <= 1'b1;
                  spc318_inst_done         <= `ARIANE_CORE318.piton_pc_vld;
                  spc318_phy_pc_w          <= `ARIANE_CORE318.piton_pc;
                end
            end
    

            assign spc319_thread_id = 2'b00;
            assign spc319_rtl_pc = spc319_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(319*4)]   <= 1'b0;
                  active_thread[(319*4)+1] <= 1'b0;
                  active_thread[(319*4)+2] <= 1'b0;
                  active_thread[(319*4)+3] <= 1'b0;
                  spc319_inst_done         <= 0;
                  spc319_phy_pc_w          <= 0;
                end else begin
                  active_thread[(319*4)]   <= 1'b1;
                  active_thread[(319*4)+1] <= 1'b1;
                  active_thread[(319*4)+2] <= 1'b1;
                  active_thread[(319*4)+3] <= 1'b1;
                  spc319_inst_done         <= `ARIANE_CORE319.piton_pc_vld;
                  spc319_phy_pc_w          <= `ARIANE_CORE319.piton_pc;
                end
            end
    

            assign spc320_thread_id = 2'b00;
            assign spc320_rtl_pc = spc320_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(320*4)]   <= 1'b0;
                  active_thread[(320*4)+1] <= 1'b0;
                  active_thread[(320*4)+2] <= 1'b0;
                  active_thread[(320*4)+3] <= 1'b0;
                  spc320_inst_done         <= 0;
                  spc320_phy_pc_w          <= 0;
                end else begin
                  active_thread[(320*4)]   <= 1'b1;
                  active_thread[(320*4)+1] <= 1'b1;
                  active_thread[(320*4)+2] <= 1'b1;
                  active_thread[(320*4)+3] <= 1'b1;
                  spc320_inst_done         <= `ARIANE_CORE320.piton_pc_vld;
                  spc320_phy_pc_w          <= `ARIANE_CORE320.piton_pc;
                end
            end
    

            assign spc321_thread_id = 2'b00;
            assign spc321_rtl_pc = spc321_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(321*4)]   <= 1'b0;
                  active_thread[(321*4)+1] <= 1'b0;
                  active_thread[(321*4)+2] <= 1'b0;
                  active_thread[(321*4)+3] <= 1'b0;
                  spc321_inst_done         <= 0;
                  spc321_phy_pc_w          <= 0;
                end else begin
                  active_thread[(321*4)]   <= 1'b1;
                  active_thread[(321*4)+1] <= 1'b1;
                  active_thread[(321*4)+2] <= 1'b1;
                  active_thread[(321*4)+3] <= 1'b1;
                  spc321_inst_done         <= `ARIANE_CORE321.piton_pc_vld;
                  spc321_phy_pc_w          <= `ARIANE_CORE321.piton_pc;
                end
            end
    

            assign spc322_thread_id = 2'b00;
            assign spc322_rtl_pc = spc322_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(322*4)]   <= 1'b0;
                  active_thread[(322*4)+1] <= 1'b0;
                  active_thread[(322*4)+2] <= 1'b0;
                  active_thread[(322*4)+3] <= 1'b0;
                  spc322_inst_done         <= 0;
                  spc322_phy_pc_w          <= 0;
                end else begin
                  active_thread[(322*4)]   <= 1'b1;
                  active_thread[(322*4)+1] <= 1'b1;
                  active_thread[(322*4)+2] <= 1'b1;
                  active_thread[(322*4)+3] <= 1'b1;
                  spc322_inst_done         <= `ARIANE_CORE322.piton_pc_vld;
                  spc322_phy_pc_w          <= `ARIANE_CORE322.piton_pc;
                end
            end
    

            assign spc323_thread_id = 2'b00;
            assign spc323_rtl_pc = spc323_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(323*4)]   <= 1'b0;
                  active_thread[(323*4)+1] <= 1'b0;
                  active_thread[(323*4)+2] <= 1'b0;
                  active_thread[(323*4)+3] <= 1'b0;
                  spc323_inst_done         <= 0;
                  spc323_phy_pc_w          <= 0;
                end else begin
                  active_thread[(323*4)]   <= 1'b1;
                  active_thread[(323*4)+1] <= 1'b1;
                  active_thread[(323*4)+2] <= 1'b1;
                  active_thread[(323*4)+3] <= 1'b1;
                  spc323_inst_done         <= `ARIANE_CORE323.piton_pc_vld;
                  spc323_phy_pc_w          <= `ARIANE_CORE323.piton_pc;
                end
            end
    

            assign spc324_thread_id = 2'b00;
            assign spc324_rtl_pc = spc324_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(324*4)]   <= 1'b0;
                  active_thread[(324*4)+1] <= 1'b0;
                  active_thread[(324*4)+2] <= 1'b0;
                  active_thread[(324*4)+3] <= 1'b0;
                  spc324_inst_done         <= 0;
                  spc324_phy_pc_w          <= 0;
                end else begin
                  active_thread[(324*4)]   <= 1'b1;
                  active_thread[(324*4)+1] <= 1'b1;
                  active_thread[(324*4)+2] <= 1'b1;
                  active_thread[(324*4)+3] <= 1'b1;
                  spc324_inst_done         <= `ARIANE_CORE324.piton_pc_vld;
                  spc324_phy_pc_w          <= `ARIANE_CORE324.piton_pc;
                end
            end
    

            assign spc325_thread_id = 2'b00;
            assign spc325_rtl_pc = spc325_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(325*4)]   <= 1'b0;
                  active_thread[(325*4)+1] <= 1'b0;
                  active_thread[(325*4)+2] <= 1'b0;
                  active_thread[(325*4)+3] <= 1'b0;
                  spc325_inst_done         <= 0;
                  spc325_phy_pc_w          <= 0;
                end else begin
                  active_thread[(325*4)]   <= 1'b1;
                  active_thread[(325*4)+1] <= 1'b1;
                  active_thread[(325*4)+2] <= 1'b1;
                  active_thread[(325*4)+3] <= 1'b1;
                  spc325_inst_done         <= `ARIANE_CORE325.piton_pc_vld;
                  spc325_phy_pc_w          <= `ARIANE_CORE325.piton_pc;
                end
            end
    

            assign spc326_thread_id = 2'b00;
            assign spc326_rtl_pc = spc326_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(326*4)]   <= 1'b0;
                  active_thread[(326*4)+1] <= 1'b0;
                  active_thread[(326*4)+2] <= 1'b0;
                  active_thread[(326*4)+3] <= 1'b0;
                  spc326_inst_done         <= 0;
                  spc326_phy_pc_w          <= 0;
                end else begin
                  active_thread[(326*4)]   <= 1'b1;
                  active_thread[(326*4)+1] <= 1'b1;
                  active_thread[(326*4)+2] <= 1'b1;
                  active_thread[(326*4)+3] <= 1'b1;
                  spc326_inst_done         <= `ARIANE_CORE326.piton_pc_vld;
                  spc326_phy_pc_w          <= `ARIANE_CORE326.piton_pc;
                end
            end
    

            assign spc327_thread_id = 2'b00;
            assign spc327_rtl_pc = spc327_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(327*4)]   <= 1'b0;
                  active_thread[(327*4)+1] <= 1'b0;
                  active_thread[(327*4)+2] <= 1'b0;
                  active_thread[(327*4)+3] <= 1'b0;
                  spc327_inst_done         <= 0;
                  spc327_phy_pc_w          <= 0;
                end else begin
                  active_thread[(327*4)]   <= 1'b1;
                  active_thread[(327*4)+1] <= 1'b1;
                  active_thread[(327*4)+2] <= 1'b1;
                  active_thread[(327*4)+3] <= 1'b1;
                  spc327_inst_done         <= `ARIANE_CORE327.piton_pc_vld;
                  spc327_phy_pc_w          <= `ARIANE_CORE327.piton_pc;
                end
            end
    

            assign spc328_thread_id = 2'b00;
            assign spc328_rtl_pc = spc328_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(328*4)]   <= 1'b0;
                  active_thread[(328*4)+1] <= 1'b0;
                  active_thread[(328*4)+2] <= 1'b0;
                  active_thread[(328*4)+3] <= 1'b0;
                  spc328_inst_done         <= 0;
                  spc328_phy_pc_w          <= 0;
                end else begin
                  active_thread[(328*4)]   <= 1'b1;
                  active_thread[(328*4)+1] <= 1'b1;
                  active_thread[(328*4)+2] <= 1'b1;
                  active_thread[(328*4)+3] <= 1'b1;
                  spc328_inst_done         <= `ARIANE_CORE328.piton_pc_vld;
                  spc328_phy_pc_w          <= `ARIANE_CORE328.piton_pc;
                end
            end
    

            assign spc329_thread_id = 2'b00;
            assign spc329_rtl_pc = spc329_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(329*4)]   <= 1'b0;
                  active_thread[(329*4)+1] <= 1'b0;
                  active_thread[(329*4)+2] <= 1'b0;
                  active_thread[(329*4)+3] <= 1'b0;
                  spc329_inst_done         <= 0;
                  spc329_phy_pc_w          <= 0;
                end else begin
                  active_thread[(329*4)]   <= 1'b1;
                  active_thread[(329*4)+1] <= 1'b1;
                  active_thread[(329*4)+2] <= 1'b1;
                  active_thread[(329*4)+3] <= 1'b1;
                  spc329_inst_done         <= `ARIANE_CORE329.piton_pc_vld;
                  spc329_phy_pc_w          <= `ARIANE_CORE329.piton_pc;
                end
            end
    

            assign spc330_thread_id = 2'b00;
            assign spc330_rtl_pc = spc330_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(330*4)]   <= 1'b0;
                  active_thread[(330*4)+1] <= 1'b0;
                  active_thread[(330*4)+2] <= 1'b0;
                  active_thread[(330*4)+3] <= 1'b0;
                  spc330_inst_done         <= 0;
                  spc330_phy_pc_w          <= 0;
                end else begin
                  active_thread[(330*4)]   <= 1'b1;
                  active_thread[(330*4)+1] <= 1'b1;
                  active_thread[(330*4)+2] <= 1'b1;
                  active_thread[(330*4)+3] <= 1'b1;
                  spc330_inst_done         <= `ARIANE_CORE330.piton_pc_vld;
                  spc330_phy_pc_w          <= `ARIANE_CORE330.piton_pc;
                end
            end
    

            assign spc331_thread_id = 2'b00;
            assign spc331_rtl_pc = spc331_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(331*4)]   <= 1'b0;
                  active_thread[(331*4)+1] <= 1'b0;
                  active_thread[(331*4)+2] <= 1'b0;
                  active_thread[(331*4)+3] <= 1'b0;
                  spc331_inst_done         <= 0;
                  spc331_phy_pc_w          <= 0;
                end else begin
                  active_thread[(331*4)]   <= 1'b1;
                  active_thread[(331*4)+1] <= 1'b1;
                  active_thread[(331*4)+2] <= 1'b1;
                  active_thread[(331*4)+3] <= 1'b1;
                  spc331_inst_done         <= `ARIANE_CORE331.piton_pc_vld;
                  spc331_phy_pc_w          <= `ARIANE_CORE331.piton_pc;
                end
            end
    

            assign spc332_thread_id = 2'b00;
            assign spc332_rtl_pc = spc332_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(332*4)]   <= 1'b0;
                  active_thread[(332*4)+1] <= 1'b0;
                  active_thread[(332*4)+2] <= 1'b0;
                  active_thread[(332*4)+3] <= 1'b0;
                  spc332_inst_done         <= 0;
                  spc332_phy_pc_w          <= 0;
                end else begin
                  active_thread[(332*4)]   <= 1'b1;
                  active_thread[(332*4)+1] <= 1'b1;
                  active_thread[(332*4)+2] <= 1'b1;
                  active_thread[(332*4)+3] <= 1'b1;
                  spc332_inst_done         <= `ARIANE_CORE332.piton_pc_vld;
                  spc332_phy_pc_w          <= `ARIANE_CORE332.piton_pc;
                end
            end
    

            assign spc333_thread_id = 2'b00;
            assign spc333_rtl_pc = spc333_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(333*4)]   <= 1'b0;
                  active_thread[(333*4)+1] <= 1'b0;
                  active_thread[(333*4)+2] <= 1'b0;
                  active_thread[(333*4)+3] <= 1'b0;
                  spc333_inst_done         <= 0;
                  spc333_phy_pc_w          <= 0;
                end else begin
                  active_thread[(333*4)]   <= 1'b1;
                  active_thread[(333*4)+1] <= 1'b1;
                  active_thread[(333*4)+2] <= 1'b1;
                  active_thread[(333*4)+3] <= 1'b1;
                  spc333_inst_done         <= `ARIANE_CORE333.piton_pc_vld;
                  spc333_phy_pc_w          <= `ARIANE_CORE333.piton_pc;
                end
            end
    

            assign spc334_thread_id = 2'b00;
            assign spc334_rtl_pc = spc334_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(334*4)]   <= 1'b0;
                  active_thread[(334*4)+1] <= 1'b0;
                  active_thread[(334*4)+2] <= 1'b0;
                  active_thread[(334*4)+3] <= 1'b0;
                  spc334_inst_done         <= 0;
                  spc334_phy_pc_w          <= 0;
                end else begin
                  active_thread[(334*4)]   <= 1'b1;
                  active_thread[(334*4)+1] <= 1'b1;
                  active_thread[(334*4)+2] <= 1'b1;
                  active_thread[(334*4)+3] <= 1'b1;
                  spc334_inst_done         <= `ARIANE_CORE334.piton_pc_vld;
                  spc334_phy_pc_w          <= `ARIANE_CORE334.piton_pc;
                end
            end
    

            assign spc335_thread_id = 2'b00;
            assign spc335_rtl_pc = spc335_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(335*4)]   <= 1'b0;
                  active_thread[(335*4)+1] <= 1'b0;
                  active_thread[(335*4)+2] <= 1'b0;
                  active_thread[(335*4)+3] <= 1'b0;
                  spc335_inst_done         <= 0;
                  spc335_phy_pc_w          <= 0;
                end else begin
                  active_thread[(335*4)]   <= 1'b1;
                  active_thread[(335*4)+1] <= 1'b1;
                  active_thread[(335*4)+2] <= 1'b1;
                  active_thread[(335*4)+3] <= 1'b1;
                  spc335_inst_done         <= `ARIANE_CORE335.piton_pc_vld;
                  spc335_phy_pc_w          <= `ARIANE_CORE335.piton_pc;
                end
            end
    

            assign spc336_thread_id = 2'b00;
            assign spc336_rtl_pc = spc336_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(336*4)]   <= 1'b0;
                  active_thread[(336*4)+1] <= 1'b0;
                  active_thread[(336*4)+2] <= 1'b0;
                  active_thread[(336*4)+3] <= 1'b0;
                  spc336_inst_done         <= 0;
                  spc336_phy_pc_w          <= 0;
                end else begin
                  active_thread[(336*4)]   <= 1'b1;
                  active_thread[(336*4)+1] <= 1'b1;
                  active_thread[(336*4)+2] <= 1'b1;
                  active_thread[(336*4)+3] <= 1'b1;
                  spc336_inst_done         <= `ARIANE_CORE336.piton_pc_vld;
                  spc336_phy_pc_w          <= `ARIANE_CORE336.piton_pc;
                end
            end
    

            assign spc337_thread_id = 2'b00;
            assign spc337_rtl_pc = spc337_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(337*4)]   <= 1'b0;
                  active_thread[(337*4)+1] <= 1'b0;
                  active_thread[(337*4)+2] <= 1'b0;
                  active_thread[(337*4)+3] <= 1'b0;
                  spc337_inst_done         <= 0;
                  spc337_phy_pc_w          <= 0;
                end else begin
                  active_thread[(337*4)]   <= 1'b1;
                  active_thread[(337*4)+1] <= 1'b1;
                  active_thread[(337*4)+2] <= 1'b1;
                  active_thread[(337*4)+3] <= 1'b1;
                  spc337_inst_done         <= `ARIANE_CORE337.piton_pc_vld;
                  spc337_phy_pc_w          <= `ARIANE_CORE337.piton_pc;
                end
            end
    

            assign spc338_thread_id = 2'b00;
            assign spc338_rtl_pc = spc338_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(338*4)]   <= 1'b0;
                  active_thread[(338*4)+1] <= 1'b0;
                  active_thread[(338*4)+2] <= 1'b0;
                  active_thread[(338*4)+3] <= 1'b0;
                  spc338_inst_done         <= 0;
                  spc338_phy_pc_w          <= 0;
                end else begin
                  active_thread[(338*4)]   <= 1'b1;
                  active_thread[(338*4)+1] <= 1'b1;
                  active_thread[(338*4)+2] <= 1'b1;
                  active_thread[(338*4)+3] <= 1'b1;
                  spc338_inst_done         <= `ARIANE_CORE338.piton_pc_vld;
                  spc338_phy_pc_w          <= `ARIANE_CORE338.piton_pc;
                end
            end
    

            assign spc339_thread_id = 2'b00;
            assign spc339_rtl_pc = spc339_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(339*4)]   <= 1'b0;
                  active_thread[(339*4)+1] <= 1'b0;
                  active_thread[(339*4)+2] <= 1'b0;
                  active_thread[(339*4)+3] <= 1'b0;
                  spc339_inst_done         <= 0;
                  spc339_phy_pc_w          <= 0;
                end else begin
                  active_thread[(339*4)]   <= 1'b1;
                  active_thread[(339*4)+1] <= 1'b1;
                  active_thread[(339*4)+2] <= 1'b1;
                  active_thread[(339*4)+3] <= 1'b1;
                  spc339_inst_done         <= `ARIANE_CORE339.piton_pc_vld;
                  spc339_phy_pc_w          <= `ARIANE_CORE339.piton_pc;
                end
            end
    

            assign spc340_thread_id = 2'b00;
            assign spc340_rtl_pc = spc340_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(340*4)]   <= 1'b0;
                  active_thread[(340*4)+1] <= 1'b0;
                  active_thread[(340*4)+2] <= 1'b0;
                  active_thread[(340*4)+3] <= 1'b0;
                  spc340_inst_done         <= 0;
                  spc340_phy_pc_w          <= 0;
                end else begin
                  active_thread[(340*4)]   <= 1'b1;
                  active_thread[(340*4)+1] <= 1'b1;
                  active_thread[(340*4)+2] <= 1'b1;
                  active_thread[(340*4)+3] <= 1'b1;
                  spc340_inst_done         <= `ARIANE_CORE340.piton_pc_vld;
                  spc340_phy_pc_w          <= `ARIANE_CORE340.piton_pc;
                end
            end
    

            assign spc341_thread_id = 2'b00;
            assign spc341_rtl_pc = spc341_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(341*4)]   <= 1'b0;
                  active_thread[(341*4)+1] <= 1'b0;
                  active_thread[(341*4)+2] <= 1'b0;
                  active_thread[(341*4)+3] <= 1'b0;
                  spc341_inst_done         <= 0;
                  spc341_phy_pc_w          <= 0;
                end else begin
                  active_thread[(341*4)]   <= 1'b1;
                  active_thread[(341*4)+1] <= 1'b1;
                  active_thread[(341*4)+2] <= 1'b1;
                  active_thread[(341*4)+3] <= 1'b1;
                  spc341_inst_done         <= `ARIANE_CORE341.piton_pc_vld;
                  spc341_phy_pc_w          <= `ARIANE_CORE341.piton_pc;
                end
            end
    

            assign spc342_thread_id = 2'b00;
            assign spc342_rtl_pc = spc342_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(342*4)]   <= 1'b0;
                  active_thread[(342*4)+1] <= 1'b0;
                  active_thread[(342*4)+2] <= 1'b0;
                  active_thread[(342*4)+3] <= 1'b0;
                  spc342_inst_done         <= 0;
                  spc342_phy_pc_w          <= 0;
                end else begin
                  active_thread[(342*4)]   <= 1'b1;
                  active_thread[(342*4)+1] <= 1'b1;
                  active_thread[(342*4)+2] <= 1'b1;
                  active_thread[(342*4)+3] <= 1'b1;
                  spc342_inst_done         <= `ARIANE_CORE342.piton_pc_vld;
                  spc342_phy_pc_w          <= `ARIANE_CORE342.piton_pc;
                end
            end
    

            assign spc343_thread_id = 2'b00;
            assign spc343_rtl_pc = spc343_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(343*4)]   <= 1'b0;
                  active_thread[(343*4)+1] <= 1'b0;
                  active_thread[(343*4)+2] <= 1'b0;
                  active_thread[(343*4)+3] <= 1'b0;
                  spc343_inst_done         <= 0;
                  spc343_phy_pc_w          <= 0;
                end else begin
                  active_thread[(343*4)]   <= 1'b1;
                  active_thread[(343*4)+1] <= 1'b1;
                  active_thread[(343*4)+2] <= 1'b1;
                  active_thread[(343*4)+3] <= 1'b1;
                  spc343_inst_done         <= `ARIANE_CORE343.piton_pc_vld;
                  spc343_phy_pc_w          <= `ARIANE_CORE343.piton_pc;
                end
            end
    

            assign spc344_thread_id = 2'b00;
            assign spc344_rtl_pc = spc344_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(344*4)]   <= 1'b0;
                  active_thread[(344*4)+1] <= 1'b0;
                  active_thread[(344*4)+2] <= 1'b0;
                  active_thread[(344*4)+3] <= 1'b0;
                  spc344_inst_done         <= 0;
                  spc344_phy_pc_w          <= 0;
                end else begin
                  active_thread[(344*4)]   <= 1'b1;
                  active_thread[(344*4)+1] <= 1'b1;
                  active_thread[(344*4)+2] <= 1'b1;
                  active_thread[(344*4)+3] <= 1'b1;
                  spc344_inst_done         <= `ARIANE_CORE344.piton_pc_vld;
                  spc344_phy_pc_w          <= `ARIANE_CORE344.piton_pc;
                end
            end
    

            assign spc345_thread_id = 2'b00;
            assign spc345_rtl_pc = spc345_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(345*4)]   <= 1'b0;
                  active_thread[(345*4)+1] <= 1'b0;
                  active_thread[(345*4)+2] <= 1'b0;
                  active_thread[(345*4)+3] <= 1'b0;
                  spc345_inst_done         <= 0;
                  spc345_phy_pc_w          <= 0;
                end else begin
                  active_thread[(345*4)]   <= 1'b1;
                  active_thread[(345*4)+1] <= 1'b1;
                  active_thread[(345*4)+2] <= 1'b1;
                  active_thread[(345*4)+3] <= 1'b1;
                  spc345_inst_done         <= `ARIANE_CORE345.piton_pc_vld;
                  spc345_phy_pc_w          <= `ARIANE_CORE345.piton_pc;
                end
            end
    

            assign spc346_thread_id = 2'b00;
            assign spc346_rtl_pc = spc346_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(346*4)]   <= 1'b0;
                  active_thread[(346*4)+1] <= 1'b0;
                  active_thread[(346*4)+2] <= 1'b0;
                  active_thread[(346*4)+3] <= 1'b0;
                  spc346_inst_done         <= 0;
                  spc346_phy_pc_w          <= 0;
                end else begin
                  active_thread[(346*4)]   <= 1'b1;
                  active_thread[(346*4)+1] <= 1'b1;
                  active_thread[(346*4)+2] <= 1'b1;
                  active_thread[(346*4)+3] <= 1'b1;
                  spc346_inst_done         <= `ARIANE_CORE346.piton_pc_vld;
                  spc346_phy_pc_w          <= `ARIANE_CORE346.piton_pc;
                end
            end
    

            assign spc347_thread_id = 2'b00;
            assign spc347_rtl_pc = spc347_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(347*4)]   <= 1'b0;
                  active_thread[(347*4)+1] <= 1'b0;
                  active_thread[(347*4)+2] <= 1'b0;
                  active_thread[(347*4)+3] <= 1'b0;
                  spc347_inst_done         <= 0;
                  spc347_phy_pc_w          <= 0;
                end else begin
                  active_thread[(347*4)]   <= 1'b1;
                  active_thread[(347*4)+1] <= 1'b1;
                  active_thread[(347*4)+2] <= 1'b1;
                  active_thread[(347*4)+3] <= 1'b1;
                  spc347_inst_done         <= `ARIANE_CORE347.piton_pc_vld;
                  spc347_phy_pc_w          <= `ARIANE_CORE347.piton_pc;
                end
            end
    

            assign spc348_thread_id = 2'b00;
            assign spc348_rtl_pc = spc348_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(348*4)]   <= 1'b0;
                  active_thread[(348*4)+1] <= 1'b0;
                  active_thread[(348*4)+2] <= 1'b0;
                  active_thread[(348*4)+3] <= 1'b0;
                  spc348_inst_done         <= 0;
                  spc348_phy_pc_w          <= 0;
                end else begin
                  active_thread[(348*4)]   <= 1'b1;
                  active_thread[(348*4)+1] <= 1'b1;
                  active_thread[(348*4)+2] <= 1'b1;
                  active_thread[(348*4)+3] <= 1'b1;
                  spc348_inst_done         <= `ARIANE_CORE348.piton_pc_vld;
                  spc348_phy_pc_w          <= `ARIANE_CORE348.piton_pc;
                end
            end
    

            assign spc349_thread_id = 2'b00;
            assign spc349_rtl_pc = spc349_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(349*4)]   <= 1'b0;
                  active_thread[(349*4)+1] <= 1'b0;
                  active_thread[(349*4)+2] <= 1'b0;
                  active_thread[(349*4)+3] <= 1'b0;
                  spc349_inst_done         <= 0;
                  spc349_phy_pc_w          <= 0;
                end else begin
                  active_thread[(349*4)]   <= 1'b1;
                  active_thread[(349*4)+1] <= 1'b1;
                  active_thread[(349*4)+2] <= 1'b1;
                  active_thread[(349*4)+3] <= 1'b1;
                  spc349_inst_done         <= `ARIANE_CORE349.piton_pc_vld;
                  spc349_phy_pc_w          <= `ARIANE_CORE349.piton_pc;
                end
            end
    

            assign spc350_thread_id = 2'b00;
            assign spc350_rtl_pc = spc350_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(350*4)]   <= 1'b0;
                  active_thread[(350*4)+1] <= 1'b0;
                  active_thread[(350*4)+2] <= 1'b0;
                  active_thread[(350*4)+3] <= 1'b0;
                  spc350_inst_done         <= 0;
                  spc350_phy_pc_w          <= 0;
                end else begin
                  active_thread[(350*4)]   <= 1'b1;
                  active_thread[(350*4)+1] <= 1'b1;
                  active_thread[(350*4)+2] <= 1'b1;
                  active_thread[(350*4)+3] <= 1'b1;
                  spc350_inst_done         <= `ARIANE_CORE350.piton_pc_vld;
                  spc350_phy_pc_w          <= `ARIANE_CORE350.piton_pc;
                end
            end
    

            assign spc351_thread_id = 2'b00;
            assign spc351_rtl_pc = spc351_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(351*4)]   <= 1'b0;
                  active_thread[(351*4)+1] <= 1'b0;
                  active_thread[(351*4)+2] <= 1'b0;
                  active_thread[(351*4)+3] <= 1'b0;
                  spc351_inst_done         <= 0;
                  spc351_phy_pc_w          <= 0;
                end else begin
                  active_thread[(351*4)]   <= 1'b1;
                  active_thread[(351*4)+1] <= 1'b1;
                  active_thread[(351*4)+2] <= 1'b1;
                  active_thread[(351*4)+3] <= 1'b1;
                  spc351_inst_done         <= `ARIANE_CORE351.piton_pc_vld;
                  spc351_phy_pc_w          <= `ARIANE_CORE351.piton_pc;
                end
            end
    

            assign spc352_thread_id = 2'b00;
            assign spc352_rtl_pc = spc352_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(352*4)]   <= 1'b0;
                  active_thread[(352*4)+1] <= 1'b0;
                  active_thread[(352*4)+2] <= 1'b0;
                  active_thread[(352*4)+3] <= 1'b0;
                  spc352_inst_done         <= 0;
                  spc352_phy_pc_w          <= 0;
                end else begin
                  active_thread[(352*4)]   <= 1'b1;
                  active_thread[(352*4)+1] <= 1'b1;
                  active_thread[(352*4)+2] <= 1'b1;
                  active_thread[(352*4)+3] <= 1'b1;
                  spc352_inst_done         <= `ARIANE_CORE352.piton_pc_vld;
                  spc352_phy_pc_w          <= `ARIANE_CORE352.piton_pc;
                end
            end
    

            assign spc353_thread_id = 2'b00;
            assign spc353_rtl_pc = spc353_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(353*4)]   <= 1'b0;
                  active_thread[(353*4)+1] <= 1'b0;
                  active_thread[(353*4)+2] <= 1'b0;
                  active_thread[(353*4)+3] <= 1'b0;
                  spc353_inst_done         <= 0;
                  spc353_phy_pc_w          <= 0;
                end else begin
                  active_thread[(353*4)]   <= 1'b1;
                  active_thread[(353*4)+1] <= 1'b1;
                  active_thread[(353*4)+2] <= 1'b1;
                  active_thread[(353*4)+3] <= 1'b1;
                  spc353_inst_done         <= `ARIANE_CORE353.piton_pc_vld;
                  spc353_phy_pc_w          <= `ARIANE_CORE353.piton_pc;
                end
            end
    

            assign spc354_thread_id = 2'b00;
            assign spc354_rtl_pc = spc354_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(354*4)]   <= 1'b0;
                  active_thread[(354*4)+1] <= 1'b0;
                  active_thread[(354*4)+2] <= 1'b0;
                  active_thread[(354*4)+3] <= 1'b0;
                  spc354_inst_done         <= 0;
                  spc354_phy_pc_w          <= 0;
                end else begin
                  active_thread[(354*4)]   <= 1'b1;
                  active_thread[(354*4)+1] <= 1'b1;
                  active_thread[(354*4)+2] <= 1'b1;
                  active_thread[(354*4)+3] <= 1'b1;
                  spc354_inst_done         <= `ARIANE_CORE354.piton_pc_vld;
                  spc354_phy_pc_w          <= `ARIANE_CORE354.piton_pc;
                end
            end
    

            assign spc355_thread_id = 2'b00;
            assign spc355_rtl_pc = spc355_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(355*4)]   <= 1'b0;
                  active_thread[(355*4)+1] <= 1'b0;
                  active_thread[(355*4)+2] <= 1'b0;
                  active_thread[(355*4)+3] <= 1'b0;
                  spc355_inst_done         <= 0;
                  spc355_phy_pc_w          <= 0;
                end else begin
                  active_thread[(355*4)]   <= 1'b1;
                  active_thread[(355*4)+1] <= 1'b1;
                  active_thread[(355*4)+2] <= 1'b1;
                  active_thread[(355*4)+3] <= 1'b1;
                  spc355_inst_done         <= `ARIANE_CORE355.piton_pc_vld;
                  spc355_phy_pc_w          <= `ARIANE_CORE355.piton_pc;
                end
            end
    

            assign spc356_thread_id = 2'b00;
            assign spc356_rtl_pc = spc356_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(356*4)]   <= 1'b0;
                  active_thread[(356*4)+1] <= 1'b0;
                  active_thread[(356*4)+2] <= 1'b0;
                  active_thread[(356*4)+3] <= 1'b0;
                  spc356_inst_done         <= 0;
                  spc356_phy_pc_w          <= 0;
                end else begin
                  active_thread[(356*4)]   <= 1'b1;
                  active_thread[(356*4)+1] <= 1'b1;
                  active_thread[(356*4)+2] <= 1'b1;
                  active_thread[(356*4)+3] <= 1'b1;
                  spc356_inst_done         <= `ARIANE_CORE356.piton_pc_vld;
                  spc356_phy_pc_w          <= `ARIANE_CORE356.piton_pc;
                end
            end
    

            assign spc357_thread_id = 2'b00;
            assign spc357_rtl_pc = spc357_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(357*4)]   <= 1'b0;
                  active_thread[(357*4)+1] <= 1'b0;
                  active_thread[(357*4)+2] <= 1'b0;
                  active_thread[(357*4)+3] <= 1'b0;
                  spc357_inst_done         <= 0;
                  spc357_phy_pc_w          <= 0;
                end else begin
                  active_thread[(357*4)]   <= 1'b1;
                  active_thread[(357*4)+1] <= 1'b1;
                  active_thread[(357*4)+2] <= 1'b1;
                  active_thread[(357*4)+3] <= 1'b1;
                  spc357_inst_done         <= `ARIANE_CORE357.piton_pc_vld;
                  spc357_phy_pc_w          <= `ARIANE_CORE357.piton_pc;
                end
            end
    

            assign spc358_thread_id = 2'b00;
            assign spc358_rtl_pc = spc358_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(358*4)]   <= 1'b0;
                  active_thread[(358*4)+1] <= 1'b0;
                  active_thread[(358*4)+2] <= 1'b0;
                  active_thread[(358*4)+3] <= 1'b0;
                  spc358_inst_done         <= 0;
                  spc358_phy_pc_w          <= 0;
                end else begin
                  active_thread[(358*4)]   <= 1'b1;
                  active_thread[(358*4)+1] <= 1'b1;
                  active_thread[(358*4)+2] <= 1'b1;
                  active_thread[(358*4)+3] <= 1'b1;
                  spc358_inst_done         <= `ARIANE_CORE358.piton_pc_vld;
                  spc358_phy_pc_w          <= `ARIANE_CORE358.piton_pc;
                end
            end
    

            assign spc359_thread_id = 2'b00;
            assign spc359_rtl_pc = spc359_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(359*4)]   <= 1'b0;
                  active_thread[(359*4)+1] <= 1'b0;
                  active_thread[(359*4)+2] <= 1'b0;
                  active_thread[(359*4)+3] <= 1'b0;
                  spc359_inst_done         <= 0;
                  spc359_phy_pc_w          <= 0;
                end else begin
                  active_thread[(359*4)]   <= 1'b1;
                  active_thread[(359*4)+1] <= 1'b1;
                  active_thread[(359*4)+2] <= 1'b1;
                  active_thread[(359*4)+3] <= 1'b1;
                  spc359_inst_done         <= `ARIANE_CORE359.piton_pc_vld;
                  spc359_phy_pc_w          <= `ARIANE_CORE359.piton_pc;
                end
            end
    

            assign spc360_thread_id = 2'b00;
            assign spc360_rtl_pc = spc360_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(360*4)]   <= 1'b0;
                  active_thread[(360*4)+1] <= 1'b0;
                  active_thread[(360*4)+2] <= 1'b0;
                  active_thread[(360*4)+3] <= 1'b0;
                  spc360_inst_done         <= 0;
                  spc360_phy_pc_w          <= 0;
                end else begin
                  active_thread[(360*4)]   <= 1'b1;
                  active_thread[(360*4)+1] <= 1'b1;
                  active_thread[(360*4)+2] <= 1'b1;
                  active_thread[(360*4)+3] <= 1'b1;
                  spc360_inst_done         <= `ARIANE_CORE360.piton_pc_vld;
                  spc360_phy_pc_w          <= `ARIANE_CORE360.piton_pc;
                end
            end
    

            assign spc361_thread_id = 2'b00;
            assign spc361_rtl_pc = spc361_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(361*4)]   <= 1'b0;
                  active_thread[(361*4)+1] <= 1'b0;
                  active_thread[(361*4)+2] <= 1'b0;
                  active_thread[(361*4)+3] <= 1'b0;
                  spc361_inst_done         <= 0;
                  spc361_phy_pc_w          <= 0;
                end else begin
                  active_thread[(361*4)]   <= 1'b1;
                  active_thread[(361*4)+1] <= 1'b1;
                  active_thread[(361*4)+2] <= 1'b1;
                  active_thread[(361*4)+3] <= 1'b1;
                  spc361_inst_done         <= `ARIANE_CORE361.piton_pc_vld;
                  spc361_phy_pc_w          <= `ARIANE_CORE361.piton_pc;
                end
            end
    

            assign spc362_thread_id = 2'b00;
            assign spc362_rtl_pc = spc362_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(362*4)]   <= 1'b0;
                  active_thread[(362*4)+1] <= 1'b0;
                  active_thread[(362*4)+2] <= 1'b0;
                  active_thread[(362*4)+3] <= 1'b0;
                  spc362_inst_done         <= 0;
                  spc362_phy_pc_w          <= 0;
                end else begin
                  active_thread[(362*4)]   <= 1'b1;
                  active_thread[(362*4)+1] <= 1'b1;
                  active_thread[(362*4)+2] <= 1'b1;
                  active_thread[(362*4)+3] <= 1'b1;
                  spc362_inst_done         <= `ARIANE_CORE362.piton_pc_vld;
                  spc362_phy_pc_w          <= `ARIANE_CORE362.piton_pc;
                end
            end
    

            assign spc363_thread_id = 2'b00;
            assign spc363_rtl_pc = spc363_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(363*4)]   <= 1'b0;
                  active_thread[(363*4)+1] <= 1'b0;
                  active_thread[(363*4)+2] <= 1'b0;
                  active_thread[(363*4)+3] <= 1'b0;
                  spc363_inst_done         <= 0;
                  spc363_phy_pc_w          <= 0;
                end else begin
                  active_thread[(363*4)]   <= 1'b1;
                  active_thread[(363*4)+1] <= 1'b1;
                  active_thread[(363*4)+2] <= 1'b1;
                  active_thread[(363*4)+3] <= 1'b1;
                  spc363_inst_done         <= `ARIANE_CORE363.piton_pc_vld;
                  spc363_phy_pc_w          <= `ARIANE_CORE363.piton_pc;
                end
            end
    

            assign spc364_thread_id = 2'b00;
            assign spc364_rtl_pc = spc364_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(364*4)]   <= 1'b0;
                  active_thread[(364*4)+1] <= 1'b0;
                  active_thread[(364*4)+2] <= 1'b0;
                  active_thread[(364*4)+3] <= 1'b0;
                  spc364_inst_done         <= 0;
                  spc364_phy_pc_w          <= 0;
                end else begin
                  active_thread[(364*4)]   <= 1'b1;
                  active_thread[(364*4)+1] <= 1'b1;
                  active_thread[(364*4)+2] <= 1'b1;
                  active_thread[(364*4)+3] <= 1'b1;
                  spc364_inst_done         <= `ARIANE_CORE364.piton_pc_vld;
                  spc364_phy_pc_w          <= `ARIANE_CORE364.piton_pc;
                end
            end
    

            assign spc365_thread_id = 2'b00;
            assign spc365_rtl_pc = spc365_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(365*4)]   <= 1'b0;
                  active_thread[(365*4)+1] <= 1'b0;
                  active_thread[(365*4)+2] <= 1'b0;
                  active_thread[(365*4)+3] <= 1'b0;
                  spc365_inst_done         <= 0;
                  spc365_phy_pc_w          <= 0;
                end else begin
                  active_thread[(365*4)]   <= 1'b1;
                  active_thread[(365*4)+1] <= 1'b1;
                  active_thread[(365*4)+2] <= 1'b1;
                  active_thread[(365*4)+3] <= 1'b1;
                  spc365_inst_done         <= `ARIANE_CORE365.piton_pc_vld;
                  spc365_phy_pc_w          <= `ARIANE_CORE365.piton_pc;
                end
            end
    

            assign spc366_thread_id = 2'b00;
            assign spc366_rtl_pc = spc366_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(366*4)]   <= 1'b0;
                  active_thread[(366*4)+1] <= 1'b0;
                  active_thread[(366*4)+2] <= 1'b0;
                  active_thread[(366*4)+3] <= 1'b0;
                  spc366_inst_done         <= 0;
                  spc366_phy_pc_w          <= 0;
                end else begin
                  active_thread[(366*4)]   <= 1'b1;
                  active_thread[(366*4)+1] <= 1'b1;
                  active_thread[(366*4)+2] <= 1'b1;
                  active_thread[(366*4)+3] <= 1'b1;
                  spc366_inst_done         <= `ARIANE_CORE366.piton_pc_vld;
                  spc366_phy_pc_w          <= `ARIANE_CORE366.piton_pc;
                end
            end
    

            assign spc367_thread_id = 2'b00;
            assign spc367_rtl_pc = spc367_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(367*4)]   <= 1'b0;
                  active_thread[(367*4)+1] <= 1'b0;
                  active_thread[(367*4)+2] <= 1'b0;
                  active_thread[(367*4)+3] <= 1'b0;
                  spc367_inst_done         <= 0;
                  spc367_phy_pc_w          <= 0;
                end else begin
                  active_thread[(367*4)]   <= 1'b1;
                  active_thread[(367*4)+1] <= 1'b1;
                  active_thread[(367*4)+2] <= 1'b1;
                  active_thread[(367*4)+3] <= 1'b1;
                  spc367_inst_done         <= `ARIANE_CORE367.piton_pc_vld;
                  spc367_phy_pc_w          <= `ARIANE_CORE367.piton_pc;
                end
            end
    

            assign spc368_thread_id = 2'b00;
            assign spc368_rtl_pc = spc368_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(368*4)]   <= 1'b0;
                  active_thread[(368*4)+1] <= 1'b0;
                  active_thread[(368*4)+2] <= 1'b0;
                  active_thread[(368*4)+3] <= 1'b0;
                  spc368_inst_done         <= 0;
                  spc368_phy_pc_w          <= 0;
                end else begin
                  active_thread[(368*4)]   <= 1'b1;
                  active_thread[(368*4)+1] <= 1'b1;
                  active_thread[(368*4)+2] <= 1'b1;
                  active_thread[(368*4)+3] <= 1'b1;
                  spc368_inst_done         <= `ARIANE_CORE368.piton_pc_vld;
                  spc368_phy_pc_w          <= `ARIANE_CORE368.piton_pc;
                end
            end
    

            assign spc369_thread_id = 2'b00;
            assign spc369_rtl_pc = spc369_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(369*4)]   <= 1'b0;
                  active_thread[(369*4)+1] <= 1'b0;
                  active_thread[(369*4)+2] <= 1'b0;
                  active_thread[(369*4)+3] <= 1'b0;
                  spc369_inst_done         <= 0;
                  spc369_phy_pc_w          <= 0;
                end else begin
                  active_thread[(369*4)]   <= 1'b1;
                  active_thread[(369*4)+1] <= 1'b1;
                  active_thread[(369*4)+2] <= 1'b1;
                  active_thread[(369*4)+3] <= 1'b1;
                  spc369_inst_done         <= `ARIANE_CORE369.piton_pc_vld;
                  spc369_phy_pc_w          <= `ARIANE_CORE369.piton_pc;
                end
            end
    

            assign spc370_thread_id = 2'b00;
            assign spc370_rtl_pc = spc370_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(370*4)]   <= 1'b0;
                  active_thread[(370*4)+1] <= 1'b0;
                  active_thread[(370*4)+2] <= 1'b0;
                  active_thread[(370*4)+3] <= 1'b0;
                  spc370_inst_done         <= 0;
                  spc370_phy_pc_w          <= 0;
                end else begin
                  active_thread[(370*4)]   <= 1'b1;
                  active_thread[(370*4)+1] <= 1'b1;
                  active_thread[(370*4)+2] <= 1'b1;
                  active_thread[(370*4)+3] <= 1'b1;
                  spc370_inst_done         <= `ARIANE_CORE370.piton_pc_vld;
                  spc370_phy_pc_w          <= `ARIANE_CORE370.piton_pc;
                end
            end
    

            assign spc371_thread_id = 2'b00;
            assign spc371_rtl_pc = spc371_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(371*4)]   <= 1'b0;
                  active_thread[(371*4)+1] <= 1'b0;
                  active_thread[(371*4)+2] <= 1'b0;
                  active_thread[(371*4)+3] <= 1'b0;
                  spc371_inst_done         <= 0;
                  spc371_phy_pc_w          <= 0;
                end else begin
                  active_thread[(371*4)]   <= 1'b1;
                  active_thread[(371*4)+1] <= 1'b1;
                  active_thread[(371*4)+2] <= 1'b1;
                  active_thread[(371*4)+3] <= 1'b1;
                  spc371_inst_done         <= `ARIANE_CORE371.piton_pc_vld;
                  spc371_phy_pc_w          <= `ARIANE_CORE371.piton_pc;
                end
            end
    

            assign spc372_thread_id = 2'b00;
            assign spc372_rtl_pc = spc372_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(372*4)]   <= 1'b0;
                  active_thread[(372*4)+1] <= 1'b0;
                  active_thread[(372*4)+2] <= 1'b0;
                  active_thread[(372*4)+3] <= 1'b0;
                  spc372_inst_done         <= 0;
                  spc372_phy_pc_w          <= 0;
                end else begin
                  active_thread[(372*4)]   <= 1'b1;
                  active_thread[(372*4)+1] <= 1'b1;
                  active_thread[(372*4)+2] <= 1'b1;
                  active_thread[(372*4)+3] <= 1'b1;
                  spc372_inst_done         <= `ARIANE_CORE372.piton_pc_vld;
                  spc372_phy_pc_w          <= `ARIANE_CORE372.piton_pc;
                end
            end
    

            assign spc373_thread_id = 2'b00;
            assign spc373_rtl_pc = spc373_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(373*4)]   <= 1'b0;
                  active_thread[(373*4)+1] <= 1'b0;
                  active_thread[(373*4)+2] <= 1'b0;
                  active_thread[(373*4)+3] <= 1'b0;
                  spc373_inst_done         <= 0;
                  spc373_phy_pc_w          <= 0;
                end else begin
                  active_thread[(373*4)]   <= 1'b1;
                  active_thread[(373*4)+1] <= 1'b1;
                  active_thread[(373*4)+2] <= 1'b1;
                  active_thread[(373*4)+3] <= 1'b1;
                  spc373_inst_done         <= `ARIANE_CORE373.piton_pc_vld;
                  spc373_phy_pc_w          <= `ARIANE_CORE373.piton_pc;
                end
            end
    

            assign spc374_thread_id = 2'b00;
            assign spc374_rtl_pc = spc374_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(374*4)]   <= 1'b0;
                  active_thread[(374*4)+1] <= 1'b0;
                  active_thread[(374*4)+2] <= 1'b0;
                  active_thread[(374*4)+3] <= 1'b0;
                  spc374_inst_done         <= 0;
                  spc374_phy_pc_w          <= 0;
                end else begin
                  active_thread[(374*4)]   <= 1'b1;
                  active_thread[(374*4)+1] <= 1'b1;
                  active_thread[(374*4)+2] <= 1'b1;
                  active_thread[(374*4)+3] <= 1'b1;
                  spc374_inst_done         <= `ARIANE_CORE374.piton_pc_vld;
                  spc374_phy_pc_w          <= `ARIANE_CORE374.piton_pc;
                end
            end
    

            assign spc375_thread_id = 2'b00;
            assign spc375_rtl_pc = spc375_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(375*4)]   <= 1'b0;
                  active_thread[(375*4)+1] <= 1'b0;
                  active_thread[(375*4)+2] <= 1'b0;
                  active_thread[(375*4)+3] <= 1'b0;
                  spc375_inst_done         <= 0;
                  spc375_phy_pc_w          <= 0;
                end else begin
                  active_thread[(375*4)]   <= 1'b1;
                  active_thread[(375*4)+1] <= 1'b1;
                  active_thread[(375*4)+2] <= 1'b1;
                  active_thread[(375*4)+3] <= 1'b1;
                  spc375_inst_done         <= `ARIANE_CORE375.piton_pc_vld;
                  spc375_phy_pc_w          <= `ARIANE_CORE375.piton_pc;
                end
            end
    

            assign spc376_thread_id = 2'b00;
            assign spc376_rtl_pc = spc376_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(376*4)]   <= 1'b0;
                  active_thread[(376*4)+1] <= 1'b0;
                  active_thread[(376*4)+2] <= 1'b0;
                  active_thread[(376*4)+3] <= 1'b0;
                  spc376_inst_done         <= 0;
                  spc376_phy_pc_w          <= 0;
                end else begin
                  active_thread[(376*4)]   <= 1'b1;
                  active_thread[(376*4)+1] <= 1'b1;
                  active_thread[(376*4)+2] <= 1'b1;
                  active_thread[(376*4)+3] <= 1'b1;
                  spc376_inst_done         <= `ARIANE_CORE376.piton_pc_vld;
                  spc376_phy_pc_w          <= `ARIANE_CORE376.piton_pc;
                end
            end
    

            assign spc377_thread_id = 2'b00;
            assign spc377_rtl_pc = spc377_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(377*4)]   <= 1'b0;
                  active_thread[(377*4)+1] <= 1'b0;
                  active_thread[(377*4)+2] <= 1'b0;
                  active_thread[(377*4)+3] <= 1'b0;
                  spc377_inst_done         <= 0;
                  spc377_phy_pc_w          <= 0;
                end else begin
                  active_thread[(377*4)]   <= 1'b1;
                  active_thread[(377*4)+1] <= 1'b1;
                  active_thread[(377*4)+2] <= 1'b1;
                  active_thread[(377*4)+3] <= 1'b1;
                  spc377_inst_done         <= `ARIANE_CORE377.piton_pc_vld;
                  spc377_phy_pc_w          <= `ARIANE_CORE377.piton_pc;
                end
            end
    

            assign spc378_thread_id = 2'b00;
            assign spc378_rtl_pc = spc378_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(378*4)]   <= 1'b0;
                  active_thread[(378*4)+1] <= 1'b0;
                  active_thread[(378*4)+2] <= 1'b0;
                  active_thread[(378*4)+3] <= 1'b0;
                  spc378_inst_done         <= 0;
                  spc378_phy_pc_w          <= 0;
                end else begin
                  active_thread[(378*4)]   <= 1'b1;
                  active_thread[(378*4)+1] <= 1'b1;
                  active_thread[(378*4)+2] <= 1'b1;
                  active_thread[(378*4)+3] <= 1'b1;
                  spc378_inst_done         <= `ARIANE_CORE378.piton_pc_vld;
                  spc378_phy_pc_w          <= `ARIANE_CORE378.piton_pc;
                end
            end
    

            assign spc379_thread_id = 2'b00;
            assign spc379_rtl_pc = spc379_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(379*4)]   <= 1'b0;
                  active_thread[(379*4)+1] <= 1'b0;
                  active_thread[(379*4)+2] <= 1'b0;
                  active_thread[(379*4)+3] <= 1'b0;
                  spc379_inst_done         <= 0;
                  spc379_phy_pc_w          <= 0;
                end else begin
                  active_thread[(379*4)]   <= 1'b1;
                  active_thread[(379*4)+1] <= 1'b1;
                  active_thread[(379*4)+2] <= 1'b1;
                  active_thread[(379*4)+3] <= 1'b1;
                  spc379_inst_done         <= `ARIANE_CORE379.piton_pc_vld;
                  spc379_phy_pc_w          <= `ARIANE_CORE379.piton_pc;
                end
            end
    

            assign spc380_thread_id = 2'b00;
            assign spc380_rtl_pc = spc380_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(380*4)]   <= 1'b0;
                  active_thread[(380*4)+1] <= 1'b0;
                  active_thread[(380*4)+2] <= 1'b0;
                  active_thread[(380*4)+3] <= 1'b0;
                  spc380_inst_done         <= 0;
                  spc380_phy_pc_w          <= 0;
                end else begin
                  active_thread[(380*4)]   <= 1'b1;
                  active_thread[(380*4)+1] <= 1'b1;
                  active_thread[(380*4)+2] <= 1'b1;
                  active_thread[(380*4)+3] <= 1'b1;
                  spc380_inst_done         <= `ARIANE_CORE380.piton_pc_vld;
                  spc380_phy_pc_w          <= `ARIANE_CORE380.piton_pc;
                end
            end
    

            assign spc381_thread_id = 2'b00;
            assign spc381_rtl_pc = spc381_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(381*4)]   <= 1'b0;
                  active_thread[(381*4)+1] <= 1'b0;
                  active_thread[(381*4)+2] <= 1'b0;
                  active_thread[(381*4)+3] <= 1'b0;
                  spc381_inst_done         <= 0;
                  spc381_phy_pc_w          <= 0;
                end else begin
                  active_thread[(381*4)]   <= 1'b1;
                  active_thread[(381*4)+1] <= 1'b1;
                  active_thread[(381*4)+2] <= 1'b1;
                  active_thread[(381*4)+3] <= 1'b1;
                  spc381_inst_done         <= `ARIANE_CORE381.piton_pc_vld;
                  spc381_phy_pc_w          <= `ARIANE_CORE381.piton_pc;
                end
            end
    

            assign spc382_thread_id = 2'b00;
            assign spc382_rtl_pc = spc382_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(382*4)]   <= 1'b0;
                  active_thread[(382*4)+1] <= 1'b0;
                  active_thread[(382*4)+2] <= 1'b0;
                  active_thread[(382*4)+3] <= 1'b0;
                  spc382_inst_done         <= 0;
                  spc382_phy_pc_w          <= 0;
                end else begin
                  active_thread[(382*4)]   <= 1'b1;
                  active_thread[(382*4)+1] <= 1'b1;
                  active_thread[(382*4)+2] <= 1'b1;
                  active_thread[(382*4)+3] <= 1'b1;
                  spc382_inst_done         <= `ARIANE_CORE382.piton_pc_vld;
                  spc382_phy_pc_w          <= `ARIANE_CORE382.piton_pc;
                end
            end
    

            assign spc383_thread_id = 2'b00;
            assign spc383_rtl_pc = spc383_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(383*4)]   <= 1'b0;
                  active_thread[(383*4)+1] <= 1'b0;
                  active_thread[(383*4)+2] <= 1'b0;
                  active_thread[(383*4)+3] <= 1'b0;
                  spc383_inst_done         <= 0;
                  spc383_phy_pc_w          <= 0;
                end else begin
                  active_thread[(383*4)]   <= 1'b1;
                  active_thread[(383*4)+1] <= 1'b1;
                  active_thread[(383*4)+2] <= 1'b1;
                  active_thread[(383*4)+3] <= 1'b1;
                  spc383_inst_done         <= `ARIANE_CORE383.piton_pc_vld;
                  spc383_phy_pc_w          <= `ARIANE_CORE383.piton_pc;
                end
            end
    

            assign spc384_thread_id = 2'b00;
            assign spc384_rtl_pc = spc384_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(384*4)]   <= 1'b0;
                  active_thread[(384*4)+1] <= 1'b0;
                  active_thread[(384*4)+2] <= 1'b0;
                  active_thread[(384*4)+3] <= 1'b0;
                  spc384_inst_done         <= 0;
                  spc384_phy_pc_w          <= 0;
                end else begin
                  active_thread[(384*4)]   <= 1'b1;
                  active_thread[(384*4)+1] <= 1'b1;
                  active_thread[(384*4)+2] <= 1'b1;
                  active_thread[(384*4)+3] <= 1'b1;
                  spc384_inst_done         <= `ARIANE_CORE384.piton_pc_vld;
                  spc384_phy_pc_w          <= `ARIANE_CORE384.piton_pc;
                end
            end
    

            assign spc385_thread_id = 2'b00;
            assign spc385_rtl_pc = spc385_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(385*4)]   <= 1'b0;
                  active_thread[(385*4)+1] <= 1'b0;
                  active_thread[(385*4)+2] <= 1'b0;
                  active_thread[(385*4)+3] <= 1'b0;
                  spc385_inst_done         <= 0;
                  spc385_phy_pc_w          <= 0;
                end else begin
                  active_thread[(385*4)]   <= 1'b1;
                  active_thread[(385*4)+1] <= 1'b1;
                  active_thread[(385*4)+2] <= 1'b1;
                  active_thread[(385*4)+3] <= 1'b1;
                  spc385_inst_done         <= `ARIANE_CORE385.piton_pc_vld;
                  spc385_phy_pc_w          <= `ARIANE_CORE385.piton_pc;
                end
            end
    

            assign spc386_thread_id = 2'b00;
            assign spc386_rtl_pc = spc386_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(386*4)]   <= 1'b0;
                  active_thread[(386*4)+1] <= 1'b0;
                  active_thread[(386*4)+2] <= 1'b0;
                  active_thread[(386*4)+3] <= 1'b0;
                  spc386_inst_done         <= 0;
                  spc386_phy_pc_w          <= 0;
                end else begin
                  active_thread[(386*4)]   <= 1'b1;
                  active_thread[(386*4)+1] <= 1'b1;
                  active_thread[(386*4)+2] <= 1'b1;
                  active_thread[(386*4)+3] <= 1'b1;
                  spc386_inst_done         <= `ARIANE_CORE386.piton_pc_vld;
                  spc386_phy_pc_w          <= `ARIANE_CORE386.piton_pc;
                end
            end
    

            assign spc387_thread_id = 2'b00;
            assign spc387_rtl_pc = spc387_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(387*4)]   <= 1'b0;
                  active_thread[(387*4)+1] <= 1'b0;
                  active_thread[(387*4)+2] <= 1'b0;
                  active_thread[(387*4)+3] <= 1'b0;
                  spc387_inst_done         <= 0;
                  spc387_phy_pc_w          <= 0;
                end else begin
                  active_thread[(387*4)]   <= 1'b1;
                  active_thread[(387*4)+1] <= 1'b1;
                  active_thread[(387*4)+2] <= 1'b1;
                  active_thread[(387*4)+3] <= 1'b1;
                  spc387_inst_done         <= `ARIANE_CORE387.piton_pc_vld;
                  spc387_phy_pc_w          <= `ARIANE_CORE387.piton_pc;
                end
            end
    

            assign spc388_thread_id = 2'b00;
            assign spc388_rtl_pc = spc388_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(388*4)]   <= 1'b0;
                  active_thread[(388*4)+1] <= 1'b0;
                  active_thread[(388*4)+2] <= 1'b0;
                  active_thread[(388*4)+3] <= 1'b0;
                  spc388_inst_done         <= 0;
                  spc388_phy_pc_w          <= 0;
                end else begin
                  active_thread[(388*4)]   <= 1'b1;
                  active_thread[(388*4)+1] <= 1'b1;
                  active_thread[(388*4)+2] <= 1'b1;
                  active_thread[(388*4)+3] <= 1'b1;
                  spc388_inst_done         <= `ARIANE_CORE388.piton_pc_vld;
                  spc388_phy_pc_w          <= `ARIANE_CORE388.piton_pc;
                end
            end
    

            assign spc389_thread_id = 2'b00;
            assign spc389_rtl_pc = spc389_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(389*4)]   <= 1'b0;
                  active_thread[(389*4)+1] <= 1'b0;
                  active_thread[(389*4)+2] <= 1'b0;
                  active_thread[(389*4)+3] <= 1'b0;
                  spc389_inst_done         <= 0;
                  spc389_phy_pc_w          <= 0;
                end else begin
                  active_thread[(389*4)]   <= 1'b1;
                  active_thread[(389*4)+1] <= 1'b1;
                  active_thread[(389*4)+2] <= 1'b1;
                  active_thread[(389*4)+3] <= 1'b1;
                  spc389_inst_done         <= `ARIANE_CORE389.piton_pc_vld;
                  spc389_phy_pc_w          <= `ARIANE_CORE389.piton_pc;
                end
            end
    

            assign spc390_thread_id = 2'b00;
            assign spc390_rtl_pc = spc390_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(390*4)]   <= 1'b0;
                  active_thread[(390*4)+1] <= 1'b0;
                  active_thread[(390*4)+2] <= 1'b0;
                  active_thread[(390*4)+3] <= 1'b0;
                  spc390_inst_done         <= 0;
                  spc390_phy_pc_w          <= 0;
                end else begin
                  active_thread[(390*4)]   <= 1'b1;
                  active_thread[(390*4)+1] <= 1'b1;
                  active_thread[(390*4)+2] <= 1'b1;
                  active_thread[(390*4)+3] <= 1'b1;
                  spc390_inst_done         <= `ARIANE_CORE390.piton_pc_vld;
                  spc390_phy_pc_w          <= `ARIANE_CORE390.piton_pc;
                end
            end
    

            assign spc391_thread_id = 2'b00;
            assign spc391_rtl_pc = spc391_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(391*4)]   <= 1'b0;
                  active_thread[(391*4)+1] <= 1'b0;
                  active_thread[(391*4)+2] <= 1'b0;
                  active_thread[(391*4)+3] <= 1'b0;
                  spc391_inst_done         <= 0;
                  spc391_phy_pc_w          <= 0;
                end else begin
                  active_thread[(391*4)]   <= 1'b1;
                  active_thread[(391*4)+1] <= 1'b1;
                  active_thread[(391*4)+2] <= 1'b1;
                  active_thread[(391*4)+3] <= 1'b1;
                  spc391_inst_done         <= `ARIANE_CORE391.piton_pc_vld;
                  spc391_phy_pc_w          <= `ARIANE_CORE391.piton_pc;
                end
            end
    

            assign spc392_thread_id = 2'b00;
            assign spc392_rtl_pc = spc392_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(392*4)]   <= 1'b0;
                  active_thread[(392*4)+1] <= 1'b0;
                  active_thread[(392*4)+2] <= 1'b0;
                  active_thread[(392*4)+3] <= 1'b0;
                  spc392_inst_done         <= 0;
                  spc392_phy_pc_w          <= 0;
                end else begin
                  active_thread[(392*4)]   <= 1'b1;
                  active_thread[(392*4)+1] <= 1'b1;
                  active_thread[(392*4)+2] <= 1'b1;
                  active_thread[(392*4)+3] <= 1'b1;
                  spc392_inst_done         <= `ARIANE_CORE392.piton_pc_vld;
                  spc392_phy_pc_w          <= `ARIANE_CORE392.piton_pc;
                end
            end
    

            assign spc393_thread_id = 2'b00;
            assign spc393_rtl_pc = spc393_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(393*4)]   <= 1'b0;
                  active_thread[(393*4)+1] <= 1'b0;
                  active_thread[(393*4)+2] <= 1'b0;
                  active_thread[(393*4)+3] <= 1'b0;
                  spc393_inst_done         <= 0;
                  spc393_phy_pc_w          <= 0;
                end else begin
                  active_thread[(393*4)]   <= 1'b1;
                  active_thread[(393*4)+1] <= 1'b1;
                  active_thread[(393*4)+2] <= 1'b1;
                  active_thread[(393*4)+3] <= 1'b1;
                  spc393_inst_done         <= `ARIANE_CORE393.piton_pc_vld;
                  spc393_phy_pc_w          <= `ARIANE_CORE393.piton_pc;
                end
            end
    

            assign spc394_thread_id = 2'b00;
            assign spc394_rtl_pc = spc394_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(394*4)]   <= 1'b0;
                  active_thread[(394*4)+1] <= 1'b0;
                  active_thread[(394*4)+2] <= 1'b0;
                  active_thread[(394*4)+3] <= 1'b0;
                  spc394_inst_done         <= 0;
                  spc394_phy_pc_w          <= 0;
                end else begin
                  active_thread[(394*4)]   <= 1'b1;
                  active_thread[(394*4)+1] <= 1'b1;
                  active_thread[(394*4)+2] <= 1'b1;
                  active_thread[(394*4)+3] <= 1'b1;
                  spc394_inst_done         <= `ARIANE_CORE394.piton_pc_vld;
                  spc394_phy_pc_w          <= `ARIANE_CORE394.piton_pc;
                end
            end
    

            assign spc395_thread_id = 2'b00;
            assign spc395_rtl_pc = spc395_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(395*4)]   <= 1'b0;
                  active_thread[(395*4)+1] <= 1'b0;
                  active_thread[(395*4)+2] <= 1'b0;
                  active_thread[(395*4)+3] <= 1'b0;
                  spc395_inst_done         <= 0;
                  spc395_phy_pc_w          <= 0;
                end else begin
                  active_thread[(395*4)]   <= 1'b1;
                  active_thread[(395*4)+1] <= 1'b1;
                  active_thread[(395*4)+2] <= 1'b1;
                  active_thread[(395*4)+3] <= 1'b1;
                  spc395_inst_done         <= `ARIANE_CORE395.piton_pc_vld;
                  spc395_phy_pc_w          <= `ARIANE_CORE395.piton_pc;
                end
            end
    

            assign spc396_thread_id = 2'b00;
            assign spc396_rtl_pc = spc396_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(396*4)]   <= 1'b0;
                  active_thread[(396*4)+1] <= 1'b0;
                  active_thread[(396*4)+2] <= 1'b0;
                  active_thread[(396*4)+3] <= 1'b0;
                  spc396_inst_done         <= 0;
                  spc396_phy_pc_w          <= 0;
                end else begin
                  active_thread[(396*4)]   <= 1'b1;
                  active_thread[(396*4)+1] <= 1'b1;
                  active_thread[(396*4)+2] <= 1'b1;
                  active_thread[(396*4)+3] <= 1'b1;
                  spc396_inst_done         <= `ARIANE_CORE396.piton_pc_vld;
                  spc396_phy_pc_w          <= `ARIANE_CORE396.piton_pc;
                end
            end
    

            assign spc397_thread_id = 2'b00;
            assign spc397_rtl_pc = spc397_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(397*4)]   <= 1'b0;
                  active_thread[(397*4)+1] <= 1'b0;
                  active_thread[(397*4)+2] <= 1'b0;
                  active_thread[(397*4)+3] <= 1'b0;
                  spc397_inst_done         <= 0;
                  spc397_phy_pc_w          <= 0;
                end else begin
                  active_thread[(397*4)]   <= 1'b1;
                  active_thread[(397*4)+1] <= 1'b1;
                  active_thread[(397*4)+2] <= 1'b1;
                  active_thread[(397*4)+3] <= 1'b1;
                  spc397_inst_done         <= `ARIANE_CORE397.piton_pc_vld;
                  spc397_phy_pc_w          <= `ARIANE_CORE397.piton_pc;
                end
            end
    

            assign spc398_thread_id = 2'b00;
            assign spc398_rtl_pc = spc398_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(398*4)]   <= 1'b0;
                  active_thread[(398*4)+1] <= 1'b0;
                  active_thread[(398*4)+2] <= 1'b0;
                  active_thread[(398*4)+3] <= 1'b0;
                  spc398_inst_done         <= 0;
                  spc398_phy_pc_w          <= 0;
                end else begin
                  active_thread[(398*4)]   <= 1'b1;
                  active_thread[(398*4)+1] <= 1'b1;
                  active_thread[(398*4)+2] <= 1'b1;
                  active_thread[(398*4)+3] <= 1'b1;
                  spc398_inst_done         <= `ARIANE_CORE398.piton_pc_vld;
                  spc398_phy_pc_w          <= `ARIANE_CORE398.piton_pc;
                end
            end
    

            assign spc399_thread_id = 2'b00;
            assign spc399_rtl_pc = spc399_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(399*4)]   <= 1'b0;
                  active_thread[(399*4)+1] <= 1'b0;
                  active_thread[(399*4)+2] <= 1'b0;
                  active_thread[(399*4)+3] <= 1'b0;
                  spc399_inst_done         <= 0;
                  spc399_phy_pc_w          <= 0;
                end else begin
                  active_thread[(399*4)]   <= 1'b1;
                  active_thread[(399*4)+1] <= 1'b1;
                  active_thread[(399*4)+2] <= 1'b1;
                  active_thread[(399*4)+3] <= 1'b1;
                  spc399_inst_done         <= `ARIANE_CORE399.piton_pc_vld;
                  spc399_phy_pc_w          <= `ARIANE_CORE399.piton_pc;
                end
            end
    

            assign spc400_thread_id = 2'b00;
            assign spc400_rtl_pc = spc400_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(400*4)]   <= 1'b0;
                  active_thread[(400*4)+1] <= 1'b0;
                  active_thread[(400*4)+2] <= 1'b0;
                  active_thread[(400*4)+3] <= 1'b0;
                  spc400_inst_done         <= 0;
                  spc400_phy_pc_w          <= 0;
                end else begin
                  active_thread[(400*4)]   <= 1'b1;
                  active_thread[(400*4)+1] <= 1'b1;
                  active_thread[(400*4)+2] <= 1'b1;
                  active_thread[(400*4)+3] <= 1'b1;
                  spc400_inst_done         <= `ARIANE_CORE400.piton_pc_vld;
                  spc400_phy_pc_w          <= `ARIANE_CORE400.piton_pc;
                end
            end
    

            assign spc401_thread_id = 2'b00;
            assign spc401_rtl_pc = spc401_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(401*4)]   <= 1'b0;
                  active_thread[(401*4)+1] <= 1'b0;
                  active_thread[(401*4)+2] <= 1'b0;
                  active_thread[(401*4)+3] <= 1'b0;
                  spc401_inst_done         <= 0;
                  spc401_phy_pc_w          <= 0;
                end else begin
                  active_thread[(401*4)]   <= 1'b1;
                  active_thread[(401*4)+1] <= 1'b1;
                  active_thread[(401*4)+2] <= 1'b1;
                  active_thread[(401*4)+3] <= 1'b1;
                  spc401_inst_done         <= `ARIANE_CORE401.piton_pc_vld;
                  spc401_phy_pc_w          <= `ARIANE_CORE401.piton_pc;
                end
            end
    

            assign spc402_thread_id = 2'b00;
            assign spc402_rtl_pc = spc402_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(402*4)]   <= 1'b0;
                  active_thread[(402*4)+1] <= 1'b0;
                  active_thread[(402*4)+2] <= 1'b0;
                  active_thread[(402*4)+3] <= 1'b0;
                  spc402_inst_done         <= 0;
                  spc402_phy_pc_w          <= 0;
                end else begin
                  active_thread[(402*4)]   <= 1'b1;
                  active_thread[(402*4)+1] <= 1'b1;
                  active_thread[(402*4)+2] <= 1'b1;
                  active_thread[(402*4)+3] <= 1'b1;
                  spc402_inst_done         <= `ARIANE_CORE402.piton_pc_vld;
                  spc402_phy_pc_w          <= `ARIANE_CORE402.piton_pc;
                end
            end
    

            assign spc403_thread_id = 2'b00;
            assign spc403_rtl_pc = spc403_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(403*4)]   <= 1'b0;
                  active_thread[(403*4)+1] <= 1'b0;
                  active_thread[(403*4)+2] <= 1'b0;
                  active_thread[(403*4)+3] <= 1'b0;
                  spc403_inst_done         <= 0;
                  spc403_phy_pc_w          <= 0;
                end else begin
                  active_thread[(403*4)]   <= 1'b1;
                  active_thread[(403*4)+1] <= 1'b1;
                  active_thread[(403*4)+2] <= 1'b1;
                  active_thread[(403*4)+3] <= 1'b1;
                  spc403_inst_done         <= `ARIANE_CORE403.piton_pc_vld;
                  spc403_phy_pc_w          <= `ARIANE_CORE403.piton_pc;
                end
            end
    

            assign spc404_thread_id = 2'b00;
            assign spc404_rtl_pc = spc404_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(404*4)]   <= 1'b0;
                  active_thread[(404*4)+1] <= 1'b0;
                  active_thread[(404*4)+2] <= 1'b0;
                  active_thread[(404*4)+3] <= 1'b0;
                  spc404_inst_done         <= 0;
                  spc404_phy_pc_w          <= 0;
                end else begin
                  active_thread[(404*4)]   <= 1'b1;
                  active_thread[(404*4)+1] <= 1'b1;
                  active_thread[(404*4)+2] <= 1'b1;
                  active_thread[(404*4)+3] <= 1'b1;
                  spc404_inst_done         <= `ARIANE_CORE404.piton_pc_vld;
                  spc404_phy_pc_w          <= `ARIANE_CORE404.piton_pc;
                end
            end
    

            assign spc405_thread_id = 2'b00;
            assign spc405_rtl_pc = spc405_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(405*4)]   <= 1'b0;
                  active_thread[(405*4)+1] <= 1'b0;
                  active_thread[(405*4)+2] <= 1'b0;
                  active_thread[(405*4)+3] <= 1'b0;
                  spc405_inst_done         <= 0;
                  spc405_phy_pc_w          <= 0;
                end else begin
                  active_thread[(405*4)]   <= 1'b1;
                  active_thread[(405*4)+1] <= 1'b1;
                  active_thread[(405*4)+2] <= 1'b1;
                  active_thread[(405*4)+3] <= 1'b1;
                  spc405_inst_done         <= `ARIANE_CORE405.piton_pc_vld;
                  spc405_phy_pc_w          <= `ARIANE_CORE405.piton_pc;
                end
            end
    

            assign spc406_thread_id = 2'b00;
            assign spc406_rtl_pc = spc406_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(406*4)]   <= 1'b0;
                  active_thread[(406*4)+1] <= 1'b0;
                  active_thread[(406*4)+2] <= 1'b0;
                  active_thread[(406*4)+3] <= 1'b0;
                  spc406_inst_done         <= 0;
                  spc406_phy_pc_w          <= 0;
                end else begin
                  active_thread[(406*4)]   <= 1'b1;
                  active_thread[(406*4)+1] <= 1'b1;
                  active_thread[(406*4)+2] <= 1'b1;
                  active_thread[(406*4)+3] <= 1'b1;
                  spc406_inst_done         <= `ARIANE_CORE406.piton_pc_vld;
                  spc406_phy_pc_w          <= `ARIANE_CORE406.piton_pc;
                end
            end
    

            assign spc407_thread_id = 2'b00;
            assign spc407_rtl_pc = spc407_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(407*4)]   <= 1'b0;
                  active_thread[(407*4)+1] <= 1'b0;
                  active_thread[(407*4)+2] <= 1'b0;
                  active_thread[(407*4)+3] <= 1'b0;
                  spc407_inst_done         <= 0;
                  spc407_phy_pc_w          <= 0;
                end else begin
                  active_thread[(407*4)]   <= 1'b1;
                  active_thread[(407*4)+1] <= 1'b1;
                  active_thread[(407*4)+2] <= 1'b1;
                  active_thread[(407*4)+3] <= 1'b1;
                  spc407_inst_done         <= `ARIANE_CORE407.piton_pc_vld;
                  spc407_phy_pc_w          <= `ARIANE_CORE407.piton_pc;
                end
            end
    

            assign spc408_thread_id = 2'b00;
            assign spc408_rtl_pc = spc408_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(408*4)]   <= 1'b0;
                  active_thread[(408*4)+1] <= 1'b0;
                  active_thread[(408*4)+2] <= 1'b0;
                  active_thread[(408*4)+3] <= 1'b0;
                  spc408_inst_done         <= 0;
                  spc408_phy_pc_w          <= 0;
                end else begin
                  active_thread[(408*4)]   <= 1'b1;
                  active_thread[(408*4)+1] <= 1'b1;
                  active_thread[(408*4)+2] <= 1'b1;
                  active_thread[(408*4)+3] <= 1'b1;
                  spc408_inst_done         <= `ARIANE_CORE408.piton_pc_vld;
                  spc408_phy_pc_w          <= `ARIANE_CORE408.piton_pc;
                end
            end
    

            assign spc409_thread_id = 2'b00;
            assign spc409_rtl_pc = spc409_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(409*4)]   <= 1'b0;
                  active_thread[(409*4)+1] <= 1'b0;
                  active_thread[(409*4)+2] <= 1'b0;
                  active_thread[(409*4)+3] <= 1'b0;
                  spc409_inst_done         <= 0;
                  spc409_phy_pc_w          <= 0;
                end else begin
                  active_thread[(409*4)]   <= 1'b1;
                  active_thread[(409*4)+1] <= 1'b1;
                  active_thread[(409*4)+2] <= 1'b1;
                  active_thread[(409*4)+3] <= 1'b1;
                  spc409_inst_done         <= `ARIANE_CORE409.piton_pc_vld;
                  spc409_phy_pc_w          <= `ARIANE_CORE409.piton_pc;
                end
            end
    

            assign spc410_thread_id = 2'b00;
            assign spc410_rtl_pc = spc410_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(410*4)]   <= 1'b0;
                  active_thread[(410*4)+1] <= 1'b0;
                  active_thread[(410*4)+2] <= 1'b0;
                  active_thread[(410*4)+3] <= 1'b0;
                  spc410_inst_done         <= 0;
                  spc410_phy_pc_w          <= 0;
                end else begin
                  active_thread[(410*4)]   <= 1'b1;
                  active_thread[(410*4)+1] <= 1'b1;
                  active_thread[(410*4)+2] <= 1'b1;
                  active_thread[(410*4)+3] <= 1'b1;
                  spc410_inst_done         <= `ARIANE_CORE410.piton_pc_vld;
                  spc410_phy_pc_w          <= `ARIANE_CORE410.piton_pc;
                end
            end
    

            assign spc411_thread_id = 2'b00;
            assign spc411_rtl_pc = spc411_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(411*4)]   <= 1'b0;
                  active_thread[(411*4)+1] <= 1'b0;
                  active_thread[(411*4)+2] <= 1'b0;
                  active_thread[(411*4)+3] <= 1'b0;
                  spc411_inst_done         <= 0;
                  spc411_phy_pc_w          <= 0;
                end else begin
                  active_thread[(411*4)]   <= 1'b1;
                  active_thread[(411*4)+1] <= 1'b1;
                  active_thread[(411*4)+2] <= 1'b1;
                  active_thread[(411*4)+3] <= 1'b1;
                  spc411_inst_done         <= `ARIANE_CORE411.piton_pc_vld;
                  spc411_phy_pc_w          <= `ARIANE_CORE411.piton_pc;
                end
            end
    

            assign spc412_thread_id = 2'b00;
            assign spc412_rtl_pc = spc412_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(412*4)]   <= 1'b0;
                  active_thread[(412*4)+1] <= 1'b0;
                  active_thread[(412*4)+2] <= 1'b0;
                  active_thread[(412*4)+3] <= 1'b0;
                  spc412_inst_done         <= 0;
                  spc412_phy_pc_w          <= 0;
                end else begin
                  active_thread[(412*4)]   <= 1'b1;
                  active_thread[(412*4)+1] <= 1'b1;
                  active_thread[(412*4)+2] <= 1'b1;
                  active_thread[(412*4)+3] <= 1'b1;
                  spc412_inst_done         <= `ARIANE_CORE412.piton_pc_vld;
                  spc412_phy_pc_w          <= `ARIANE_CORE412.piton_pc;
                end
            end
    

            assign spc413_thread_id = 2'b00;
            assign spc413_rtl_pc = spc413_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(413*4)]   <= 1'b0;
                  active_thread[(413*4)+1] <= 1'b0;
                  active_thread[(413*4)+2] <= 1'b0;
                  active_thread[(413*4)+3] <= 1'b0;
                  spc413_inst_done         <= 0;
                  spc413_phy_pc_w          <= 0;
                end else begin
                  active_thread[(413*4)]   <= 1'b1;
                  active_thread[(413*4)+1] <= 1'b1;
                  active_thread[(413*4)+2] <= 1'b1;
                  active_thread[(413*4)+3] <= 1'b1;
                  spc413_inst_done         <= `ARIANE_CORE413.piton_pc_vld;
                  spc413_phy_pc_w          <= `ARIANE_CORE413.piton_pc;
                end
            end
    

            assign spc414_thread_id = 2'b00;
            assign spc414_rtl_pc = spc414_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(414*4)]   <= 1'b0;
                  active_thread[(414*4)+1] <= 1'b0;
                  active_thread[(414*4)+2] <= 1'b0;
                  active_thread[(414*4)+3] <= 1'b0;
                  spc414_inst_done         <= 0;
                  spc414_phy_pc_w          <= 0;
                end else begin
                  active_thread[(414*4)]   <= 1'b1;
                  active_thread[(414*4)+1] <= 1'b1;
                  active_thread[(414*4)+2] <= 1'b1;
                  active_thread[(414*4)+3] <= 1'b1;
                  spc414_inst_done         <= `ARIANE_CORE414.piton_pc_vld;
                  spc414_phy_pc_w          <= `ARIANE_CORE414.piton_pc;
                end
            end
    

            assign spc415_thread_id = 2'b00;
            assign spc415_rtl_pc = spc415_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(415*4)]   <= 1'b0;
                  active_thread[(415*4)+1] <= 1'b0;
                  active_thread[(415*4)+2] <= 1'b0;
                  active_thread[(415*4)+3] <= 1'b0;
                  spc415_inst_done         <= 0;
                  spc415_phy_pc_w          <= 0;
                end else begin
                  active_thread[(415*4)]   <= 1'b1;
                  active_thread[(415*4)+1] <= 1'b1;
                  active_thread[(415*4)+2] <= 1'b1;
                  active_thread[(415*4)+3] <= 1'b1;
                  spc415_inst_done         <= `ARIANE_CORE415.piton_pc_vld;
                  spc415_phy_pc_w          <= `ARIANE_CORE415.piton_pc;
                end
            end
    

            assign spc416_thread_id = 2'b00;
            assign spc416_rtl_pc = spc416_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(416*4)]   <= 1'b0;
                  active_thread[(416*4)+1] <= 1'b0;
                  active_thread[(416*4)+2] <= 1'b0;
                  active_thread[(416*4)+3] <= 1'b0;
                  spc416_inst_done         <= 0;
                  spc416_phy_pc_w          <= 0;
                end else begin
                  active_thread[(416*4)]   <= 1'b1;
                  active_thread[(416*4)+1] <= 1'b1;
                  active_thread[(416*4)+2] <= 1'b1;
                  active_thread[(416*4)+3] <= 1'b1;
                  spc416_inst_done         <= `ARIANE_CORE416.piton_pc_vld;
                  spc416_phy_pc_w          <= `ARIANE_CORE416.piton_pc;
                end
            end
    

            assign spc417_thread_id = 2'b00;
            assign spc417_rtl_pc = spc417_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(417*4)]   <= 1'b0;
                  active_thread[(417*4)+1] <= 1'b0;
                  active_thread[(417*4)+2] <= 1'b0;
                  active_thread[(417*4)+3] <= 1'b0;
                  spc417_inst_done         <= 0;
                  spc417_phy_pc_w          <= 0;
                end else begin
                  active_thread[(417*4)]   <= 1'b1;
                  active_thread[(417*4)+1] <= 1'b1;
                  active_thread[(417*4)+2] <= 1'b1;
                  active_thread[(417*4)+3] <= 1'b1;
                  spc417_inst_done         <= `ARIANE_CORE417.piton_pc_vld;
                  spc417_phy_pc_w          <= `ARIANE_CORE417.piton_pc;
                end
            end
    

            assign spc418_thread_id = 2'b00;
            assign spc418_rtl_pc = spc418_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(418*4)]   <= 1'b0;
                  active_thread[(418*4)+1] <= 1'b0;
                  active_thread[(418*4)+2] <= 1'b0;
                  active_thread[(418*4)+3] <= 1'b0;
                  spc418_inst_done         <= 0;
                  spc418_phy_pc_w          <= 0;
                end else begin
                  active_thread[(418*4)]   <= 1'b1;
                  active_thread[(418*4)+1] <= 1'b1;
                  active_thread[(418*4)+2] <= 1'b1;
                  active_thread[(418*4)+3] <= 1'b1;
                  spc418_inst_done         <= `ARIANE_CORE418.piton_pc_vld;
                  spc418_phy_pc_w          <= `ARIANE_CORE418.piton_pc;
                end
            end
    

            assign spc419_thread_id = 2'b00;
            assign spc419_rtl_pc = spc419_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(419*4)]   <= 1'b0;
                  active_thread[(419*4)+1] <= 1'b0;
                  active_thread[(419*4)+2] <= 1'b0;
                  active_thread[(419*4)+3] <= 1'b0;
                  spc419_inst_done         <= 0;
                  spc419_phy_pc_w          <= 0;
                end else begin
                  active_thread[(419*4)]   <= 1'b1;
                  active_thread[(419*4)+1] <= 1'b1;
                  active_thread[(419*4)+2] <= 1'b1;
                  active_thread[(419*4)+3] <= 1'b1;
                  spc419_inst_done         <= `ARIANE_CORE419.piton_pc_vld;
                  spc419_phy_pc_w          <= `ARIANE_CORE419.piton_pc;
                end
            end
    

            assign spc420_thread_id = 2'b00;
            assign spc420_rtl_pc = spc420_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(420*4)]   <= 1'b0;
                  active_thread[(420*4)+1] <= 1'b0;
                  active_thread[(420*4)+2] <= 1'b0;
                  active_thread[(420*4)+3] <= 1'b0;
                  spc420_inst_done         <= 0;
                  spc420_phy_pc_w          <= 0;
                end else begin
                  active_thread[(420*4)]   <= 1'b1;
                  active_thread[(420*4)+1] <= 1'b1;
                  active_thread[(420*4)+2] <= 1'b1;
                  active_thread[(420*4)+3] <= 1'b1;
                  spc420_inst_done         <= `ARIANE_CORE420.piton_pc_vld;
                  spc420_phy_pc_w          <= `ARIANE_CORE420.piton_pc;
                end
            end
    

            assign spc421_thread_id = 2'b00;
            assign spc421_rtl_pc = spc421_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(421*4)]   <= 1'b0;
                  active_thread[(421*4)+1] <= 1'b0;
                  active_thread[(421*4)+2] <= 1'b0;
                  active_thread[(421*4)+3] <= 1'b0;
                  spc421_inst_done         <= 0;
                  spc421_phy_pc_w          <= 0;
                end else begin
                  active_thread[(421*4)]   <= 1'b1;
                  active_thread[(421*4)+1] <= 1'b1;
                  active_thread[(421*4)+2] <= 1'b1;
                  active_thread[(421*4)+3] <= 1'b1;
                  spc421_inst_done         <= `ARIANE_CORE421.piton_pc_vld;
                  spc421_phy_pc_w          <= `ARIANE_CORE421.piton_pc;
                end
            end
    

            assign spc422_thread_id = 2'b00;
            assign spc422_rtl_pc = spc422_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(422*4)]   <= 1'b0;
                  active_thread[(422*4)+1] <= 1'b0;
                  active_thread[(422*4)+2] <= 1'b0;
                  active_thread[(422*4)+3] <= 1'b0;
                  spc422_inst_done         <= 0;
                  spc422_phy_pc_w          <= 0;
                end else begin
                  active_thread[(422*4)]   <= 1'b1;
                  active_thread[(422*4)+1] <= 1'b1;
                  active_thread[(422*4)+2] <= 1'b1;
                  active_thread[(422*4)+3] <= 1'b1;
                  spc422_inst_done         <= `ARIANE_CORE422.piton_pc_vld;
                  spc422_phy_pc_w          <= `ARIANE_CORE422.piton_pc;
                end
            end
    

            assign spc423_thread_id = 2'b00;
            assign spc423_rtl_pc = spc423_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(423*4)]   <= 1'b0;
                  active_thread[(423*4)+1] <= 1'b0;
                  active_thread[(423*4)+2] <= 1'b0;
                  active_thread[(423*4)+3] <= 1'b0;
                  spc423_inst_done         <= 0;
                  spc423_phy_pc_w          <= 0;
                end else begin
                  active_thread[(423*4)]   <= 1'b1;
                  active_thread[(423*4)+1] <= 1'b1;
                  active_thread[(423*4)+2] <= 1'b1;
                  active_thread[(423*4)+3] <= 1'b1;
                  spc423_inst_done         <= `ARIANE_CORE423.piton_pc_vld;
                  spc423_phy_pc_w          <= `ARIANE_CORE423.piton_pc;
                end
            end
    

            assign spc424_thread_id = 2'b00;
            assign spc424_rtl_pc = spc424_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(424*4)]   <= 1'b0;
                  active_thread[(424*4)+1] <= 1'b0;
                  active_thread[(424*4)+2] <= 1'b0;
                  active_thread[(424*4)+3] <= 1'b0;
                  spc424_inst_done         <= 0;
                  spc424_phy_pc_w          <= 0;
                end else begin
                  active_thread[(424*4)]   <= 1'b1;
                  active_thread[(424*4)+1] <= 1'b1;
                  active_thread[(424*4)+2] <= 1'b1;
                  active_thread[(424*4)+3] <= 1'b1;
                  spc424_inst_done         <= `ARIANE_CORE424.piton_pc_vld;
                  spc424_phy_pc_w          <= `ARIANE_CORE424.piton_pc;
                end
            end
    

            assign spc425_thread_id = 2'b00;
            assign spc425_rtl_pc = spc425_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(425*4)]   <= 1'b0;
                  active_thread[(425*4)+1] <= 1'b0;
                  active_thread[(425*4)+2] <= 1'b0;
                  active_thread[(425*4)+3] <= 1'b0;
                  spc425_inst_done         <= 0;
                  spc425_phy_pc_w          <= 0;
                end else begin
                  active_thread[(425*4)]   <= 1'b1;
                  active_thread[(425*4)+1] <= 1'b1;
                  active_thread[(425*4)+2] <= 1'b1;
                  active_thread[(425*4)+3] <= 1'b1;
                  spc425_inst_done         <= `ARIANE_CORE425.piton_pc_vld;
                  spc425_phy_pc_w          <= `ARIANE_CORE425.piton_pc;
                end
            end
    

            assign spc426_thread_id = 2'b00;
            assign spc426_rtl_pc = spc426_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(426*4)]   <= 1'b0;
                  active_thread[(426*4)+1] <= 1'b0;
                  active_thread[(426*4)+2] <= 1'b0;
                  active_thread[(426*4)+3] <= 1'b0;
                  spc426_inst_done         <= 0;
                  spc426_phy_pc_w          <= 0;
                end else begin
                  active_thread[(426*4)]   <= 1'b1;
                  active_thread[(426*4)+1] <= 1'b1;
                  active_thread[(426*4)+2] <= 1'b1;
                  active_thread[(426*4)+3] <= 1'b1;
                  spc426_inst_done         <= `ARIANE_CORE426.piton_pc_vld;
                  spc426_phy_pc_w          <= `ARIANE_CORE426.piton_pc;
                end
            end
    

            assign spc427_thread_id = 2'b00;
            assign spc427_rtl_pc = spc427_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(427*4)]   <= 1'b0;
                  active_thread[(427*4)+1] <= 1'b0;
                  active_thread[(427*4)+2] <= 1'b0;
                  active_thread[(427*4)+3] <= 1'b0;
                  spc427_inst_done         <= 0;
                  spc427_phy_pc_w          <= 0;
                end else begin
                  active_thread[(427*4)]   <= 1'b1;
                  active_thread[(427*4)+1] <= 1'b1;
                  active_thread[(427*4)+2] <= 1'b1;
                  active_thread[(427*4)+3] <= 1'b1;
                  spc427_inst_done         <= `ARIANE_CORE427.piton_pc_vld;
                  spc427_phy_pc_w          <= `ARIANE_CORE427.piton_pc;
                end
            end
    

            assign spc428_thread_id = 2'b00;
            assign spc428_rtl_pc = spc428_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(428*4)]   <= 1'b0;
                  active_thread[(428*4)+1] <= 1'b0;
                  active_thread[(428*4)+2] <= 1'b0;
                  active_thread[(428*4)+3] <= 1'b0;
                  spc428_inst_done         <= 0;
                  spc428_phy_pc_w          <= 0;
                end else begin
                  active_thread[(428*4)]   <= 1'b1;
                  active_thread[(428*4)+1] <= 1'b1;
                  active_thread[(428*4)+2] <= 1'b1;
                  active_thread[(428*4)+3] <= 1'b1;
                  spc428_inst_done         <= `ARIANE_CORE428.piton_pc_vld;
                  spc428_phy_pc_w          <= `ARIANE_CORE428.piton_pc;
                end
            end
    

            assign spc429_thread_id = 2'b00;
            assign spc429_rtl_pc = spc429_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(429*4)]   <= 1'b0;
                  active_thread[(429*4)+1] <= 1'b0;
                  active_thread[(429*4)+2] <= 1'b0;
                  active_thread[(429*4)+3] <= 1'b0;
                  spc429_inst_done         <= 0;
                  spc429_phy_pc_w          <= 0;
                end else begin
                  active_thread[(429*4)]   <= 1'b1;
                  active_thread[(429*4)+1] <= 1'b1;
                  active_thread[(429*4)+2] <= 1'b1;
                  active_thread[(429*4)+3] <= 1'b1;
                  spc429_inst_done         <= `ARIANE_CORE429.piton_pc_vld;
                  spc429_phy_pc_w          <= `ARIANE_CORE429.piton_pc;
                end
            end
    

            assign spc430_thread_id = 2'b00;
            assign spc430_rtl_pc = spc430_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(430*4)]   <= 1'b0;
                  active_thread[(430*4)+1] <= 1'b0;
                  active_thread[(430*4)+2] <= 1'b0;
                  active_thread[(430*4)+3] <= 1'b0;
                  spc430_inst_done         <= 0;
                  spc430_phy_pc_w          <= 0;
                end else begin
                  active_thread[(430*4)]   <= 1'b1;
                  active_thread[(430*4)+1] <= 1'b1;
                  active_thread[(430*4)+2] <= 1'b1;
                  active_thread[(430*4)+3] <= 1'b1;
                  spc430_inst_done         <= `ARIANE_CORE430.piton_pc_vld;
                  spc430_phy_pc_w          <= `ARIANE_CORE430.piton_pc;
                end
            end
    

            assign spc431_thread_id = 2'b00;
            assign spc431_rtl_pc = spc431_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(431*4)]   <= 1'b0;
                  active_thread[(431*4)+1] <= 1'b0;
                  active_thread[(431*4)+2] <= 1'b0;
                  active_thread[(431*4)+3] <= 1'b0;
                  spc431_inst_done         <= 0;
                  spc431_phy_pc_w          <= 0;
                end else begin
                  active_thread[(431*4)]   <= 1'b1;
                  active_thread[(431*4)+1] <= 1'b1;
                  active_thread[(431*4)+2] <= 1'b1;
                  active_thread[(431*4)+3] <= 1'b1;
                  spc431_inst_done         <= `ARIANE_CORE431.piton_pc_vld;
                  spc431_phy_pc_w          <= `ARIANE_CORE431.piton_pc;
                end
            end
    

            assign spc432_thread_id = 2'b00;
            assign spc432_rtl_pc = spc432_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(432*4)]   <= 1'b0;
                  active_thread[(432*4)+1] <= 1'b0;
                  active_thread[(432*4)+2] <= 1'b0;
                  active_thread[(432*4)+3] <= 1'b0;
                  spc432_inst_done         <= 0;
                  spc432_phy_pc_w          <= 0;
                end else begin
                  active_thread[(432*4)]   <= 1'b1;
                  active_thread[(432*4)+1] <= 1'b1;
                  active_thread[(432*4)+2] <= 1'b1;
                  active_thread[(432*4)+3] <= 1'b1;
                  spc432_inst_done         <= `ARIANE_CORE432.piton_pc_vld;
                  spc432_phy_pc_w          <= `ARIANE_CORE432.piton_pc;
                end
            end
    

            assign spc433_thread_id = 2'b00;
            assign spc433_rtl_pc = spc433_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(433*4)]   <= 1'b0;
                  active_thread[(433*4)+1] <= 1'b0;
                  active_thread[(433*4)+2] <= 1'b0;
                  active_thread[(433*4)+3] <= 1'b0;
                  spc433_inst_done         <= 0;
                  spc433_phy_pc_w          <= 0;
                end else begin
                  active_thread[(433*4)]   <= 1'b1;
                  active_thread[(433*4)+1] <= 1'b1;
                  active_thread[(433*4)+2] <= 1'b1;
                  active_thread[(433*4)+3] <= 1'b1;
                  spc433_inst_done         <= `ARIANE_CORE433.piton_pc_vld;
                  spc433_phy_pc_w          <= `ARIANE_CORE433.piton_pc;
                end
            end
    

            assign spc434_thread_id = 2'b00;
            assign spc434_rtl_pc = spc434_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(434*4)]   <= 1'b0;
                  active_thread[(434*4)+1] <= 1'b0;
                  active_thread[(434*4)+2] <= 1'b0;
                  active_thread[(434*4)+3] <= 1'b0;
                  spc434_inst_done         <= 0;
                  spc434_phy_pc_w          <= 0;
                end else begin
                  active_thread[(434*4)]   <= 1'b1;
                  active_thread[(434*4)+1] <= 1'b1;
                  active_thread[(434*4)+2] <= 1'b1;
                  active_thread[(434*4)+3] <= 1'b1;
                  spc434_inst_done         <= `ARIANE_CORE434.piton_pc_vld;
                  spc434_phy_pc_w          <= `ARIANE_CORE434.piton_pc;
                end
            end
    

            assign spc435_thread_id = 2'b00;
            assign spc435_rtl_pc = spc435_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(435*4)]   <= 1'b0;
                  active_thread[(435*4)+1] <= 1'b0;
                  active_thread[(435*4)+2] <= 1'b0;
                  active_thread[(435*4)+3] <= 1'b0;
                  spc435_inst_done         <= 0;
                  spc435_phy_pc_w          <= 0;
                end else begin
                  active_thread[(435*4)]   <= 1'b1;
                  active_thread[(435*4)+1] <= 1'b1;
                  active_thread[(435*4)+2] <= 1'b1;
                  active_thread[(435*4)+3] <= 1'b1;
                  spc435_inst_done         <= `ARIANE_CORE435.piton_pc_vld;
                  spc435_phy_pc_w          <= `ARIANE_CORE435.piton_pc;
                end
            end
    

            assign spc436_thread_id = 2'b00;
            assign spc436_rtl_pc = spc436_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(436*4)]   <= 1'b0;
                  active_thread[(436*4)+1] <= 1'b0;
                  active_thread[(436*4)+2] <= 1'b0;
                  active_thread[(436*4)+3] <= 1'b0;
                  spc436_inst_done         <= 0;
                  spc436_phy_pc_w          <= 0;
                end else begin
                  active_thread[(436*4)]   <= 1'b1;
                  active_thread[(436*4)+1] <= 1'b1;
                  active_thread[(436*4)+2] <= 1'b1;
                  active_thread[(436*4)+3] <= 1'b1;
                  spc436_inst_done         <= `ARIANE_CORE436.piton_pc_vld;
                  spc436_phy_pc_w          <= `ARIANE_CORE436.piton_pc;
                end
            end
    

            assign spc437_thread_id = 2'b00;
            assign spc437_rtl_pc = spc437_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(437*4)]   <= 1'b0;
                  active_thread[(437*4)+1] <= 1'b0;
                  active_thread[(437*4)+2] <= 1'b0;
                  active_thread[(437*4)+3] <= 1'b0;
                  spc437_inst_done         <= 0;
                  spc437_phy_pc_w          <= 0;
                end else begin
                  active_thread[(437*4)]   <= 1'b1;
                  active_thread[(437*4)+1] <= 1'b1;
                  active_thread[(437*4)+2] <= 1'b1;
                  active_thread[(437*4)+3] <= 1'b1;
                  spc437_inst_done         <= `ARIANE_CORE437.piton_pc_vld;
                  spc437_phy_pc_w          <= `ARIANE_CORE437.piton_pc;
                end
            end
    

            assign spc438_thread_id = 2'b00;
            assign spc438_rtl_pc = spc438_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(438*4)]   <= 1'b0;
                  active_thread[(438*4)+1] <= 1'b0;
                  active_thread[(438*4)+2] <= 1'b0;
                  active_thread[(438*4)+3] <= 1'b0;
                  spc438_inst_done         <= 0;
                  spc438_phy_pc_w          <= 0;
                end else begin
                  active_thread[(438*4)]   <= 1'b1;
                  active_thread[(438*4)+1] <= 1'b1;
                  active_thread[(438*4)+2] <= 1'b1;
                  active_thread[(438*4)+3] <= 1'b1;
                  spc438_inst_done         <= `ARIANE_CORE438.piton_pc_vld;
                  spc438_phy_pc_w          <= `ARIANE_CORE438.piton_pc;
                end
            end
    

            assign spc439_thread_id = 2'b00;
            assign spc439_rtl_pc = spc439_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(439*4)]   <= 1'b0;
                  active_thread[(439*4)+1] <= 1'b0;
                  active_thread[(439*4)+2] <= 1'b0;
                  active_thread[(439*4)+3] <= 1'b0;
                  spc439_inst_done         <= 0;
                  spc439_phy_pc_w          <= 0;
                end else begin
                  active_thread[(439*4)]   <= 1'b1;
                  active_thread[(439*4)+1] <= 1'b1;
                  active_thread[(439*4)+2] <= 1'b1;
                  active_thread[(439*4)+3] <= 1'b1;
                  spc439_inst_done         <= `ARIANE_CORE439.piton_pc_vld;
                  spc439_phy_pc_w          <= `ARIANE_CORE439.piton_pc;
                end
            end
    

            assign spc440_thread_id = 2'b00;
            assign spc440_rtl_pc = spc440_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(440*4)]   <= 1'b0;
                  active_thread[(440*4)+1] <= 1'b0;
                  active_thread[(440*4)+2] <= 1'b0;
                  active_thread[(440*4)+3] <= 1'b0;
                  spc440_inst_done         <= 0;
                  spc440_phy_pc_w          <= 0;
                end else begin
                  active_thread[(440*4)]   <= 1'b1;
                  active_thread[(440*4)+1] <= 1'b1;
                  active_thread[(440*4)+2] <= 1'b1;
                  active_thread[(440*4)+3] <= 1'b1;
                  spc440_inst_done         <= `ARIANE_CORE440.piton_pc_vld;
                  spc440_phy_pc_w          <= `ARIANE_CORE440.piton_pc;
                end
            end
    

            assign spc441_thread_id = 2'b00;
            assign spc441_rtl_pc = spc441_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(441*4)]   <= 1'b0;
                  active_thread[(441*4)+1] <= 1'b0;
                  active_thread[(441*4)+2] <= 1'b0;
                  active_thread[(441*4)+3] <= 1'b0;
                  spc441_inst_done         <= 0;
                  spc441_phy_pc_w          <= 0;
                end else begin
                  active_thread[(441*4)]   <= 1'b1;
                  active_thread[(441*4)+1] <= 1'b1;
                  active_thread[(441*4)+2] <= 1'b1;
                  active_thread[(441*4)+3] <= 1'b1;
                  spc441_inst_done         <= `ARIANE_CORE441.piton_pc_vld;
                  spc441_phy_pc_w          <= `ARIANE_CORE441.piton_pc;
                end
            end
    

            assign spc442_thread_id = 2'b00;
            assign spc442_rtl_pc = spc442_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(442*4)]   <= 1'b0;
                  active_thread[(442*4)+1] <= 1'b0;
                  active_thread[(442*4)+2] <= 1'b0;
                  active_thread[(442*4)+3] <= 1'b0;
                  spc442_inst_done         <= 0;
                  spc442_phy_pc_w          <= 0;
                end else begin
                  active_thread[(442*4)]   <= 1'b1;
                  active_thread[(442*4)+1] <= 1'b1;
                  active_thread[(442*4)+2] <= 1'b1;
                  active_thread[(442*4)+3] <= 1'b1;
                  spc442_inst_done         <= `ARIANE_CORE442.piton_pc_vld;
                  spc442_phy_pc_w          <= `ARIANE_CORE442.piton_pc;
                end
            end
    

            assign spc443_thread_id = 2'b00;
            assign spc443_rtl_pc = spc443_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(443*4)]   <= 1'b0;
                  active_thread[(443*4)+1] <= 1'b0;
                  active_thread[(443*4)+2] <= 1'b0;
                  active_thread[(443*4)+3] <= 1'b0;
                  spc443_inst_done         <= 0;
                  spc443_phy_pc_w          <= 0;
                end else begin
                  active_thread[(443*4)]   <= 1'b1;
                  active_thread[(443*4)+1] <= 1'b1;
                  active_thread[(443*4)+2] <= 1'b1;
                  active_thread[(443*4)+3] <= 1'b1;
                  spc443_inst_done         <= `ARIANE_CORE443.piton_pc_vld;
                  spc443_phy_pc_w          <= `ARIANE_CORE443.piton_pc;
                end
            end
    

            assign spc444_thread_id = 2'b00;
            assign spc444_rtl_pc = spc444_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(444*4)]   <= 1'b0;
                  active_thread[(444*4)+1] <= 1'b0;
                  active_thread[(444*4)+2] <= 1'b0;
                  active_thread[(444*4)+3] <= 1'b0;
                  spc444_inst_done         <= 0;
                  spc444_phy_pc_w          <= 0;
                end else begin
                  active_thread[(444*4)]   <= 1'b1;
                  active_thread[(444*4)+1] <= 1'b1;
                  active_thread[(444*4)+2] <= 1'b1;
                  active_thread[(444*4)+3] <= 1'b1;
                  spc444_inst_done         <= `ARIANE_CORE444.piton_pc_vld;
                  spc444_phy_pc_w          <= `ARIANE_CORE444.piton_pc;
                end
            end
    

            assign spc445_thread_id = 2'b00;
            assign spc445_rtl_pc = spc445_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(445*4)]   <= 1'b0;
                  active_thread[(445*4)+1] <= 1'b0;
                  active_thread[(445*4)+2] <= 1'b0;
                  active_thread[(445*4)+3] <= 1'b0;
                  spc445_inst_done         <= 0;
                  spc445_phy_pc_w          <= 0;
                end else begin
                  active_thread[(445*4)]   <= 1'b1;
                  active_thread[(445*4)+1] <= 1'b1;
                  active_thread[(445*4)+2] <= 1'b1;
                  active_thread[(445*4)+3] <= 1'b1;
                  spc445_inst_done         <= `ARIANE_CORE445.piton_pc_vld;
                  spc445_phy_pc_w          <= `ARIANE_CORE445.piton_pc;
                end
            end
    

            assign spc446_thread_id = 2'b00;
            assign spc446_rtl_pc = spc446_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(446*4)]   <= 1'b0;
                  active_thread[(446*4)+1] <= 1'b0;
                  active_thread[(446*4)+2] <= 1'b0;
                  active_thread[(446*4)+3] <= 1'b0;
                  spc446_inst_done         <= 0;
                  spc446_phy_pc_w          <= 0;
                end else begin
                  active_thread[(446*4)]   <= 1'b1;
                  active_thread[(446*4)+1] <= 1'b1;
                  active_thread[(446*4)+2] <= 1'b1;
                  active_thread[(446*4)+3] <= 1'b1;
                  spc446_inst_done         <= `ARIANE_CORE446.piton_pc_vld;
                  spc446_phy_pc_w          <= `ARIANE_CORE446.piton_pc;
                end
            end
    

            assign spc447_thread_id = 2'b00;
            assign spc447_rtl_pc = spc447_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(447*4)]   <= 1'b0;
                  active_thread[(447*4)+1] <= 1'b0;
                  active_thread[(447*4)+2] <= 1'b0;
                  active_thread[(447*4)+3] <= 1'b0;
                  spc447_inst_done         <= 0;
                  spc447_phy_pc_w          <= 0;
                end else begin
                  active_thread[(447*4)]   <= 1'b1;
                  active_thread[(447*4)+1] <= 1'b1;
                  active_thread[(447*4)+2] <= 1'b1;
                  active_thread[(447*4)+3] <= 1'b1;
                  spc447_inst_done         <= `ARIANE_CORE447.piton_pc_vld;
                  spc447_phy_pc_w          <= `ARIANE_CORE447.piton_pc;
                end
            end
    

            assign spc448_thread_id = 2'b00;
            assign spc448_rtl_pc = spc448_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(448*4)]   <= 1'b0;
                  active_thread[(448*4)+1] <= 1'b0;
                  active_thread[(448*4)+2] <= 1'b0;
                  active_thread[(448*4)+3] <= 1'b0;
                  spc448_inst_done         <= 0;
                  spc448_phy_pc_w          <= 0;
                end else begin
                  active_thread[(448*4)]   <= 1'b1;
                  active_thread[(448*4)+1] <= 1'b1;
                  active_thread[(448*4)+2] <= 1'b1;
                  active_thread[(448*4)+3] <= 1'b1;
                  spc448_inst_done         <= `ARIANE_CORE448.piton_pc_vld;
                  spc448_phy_pc_w          <= `ARIANE_CORE448.piton_pc;
                end
            end
    

            assign spc449_thread_id = 2'b00;
            assign spc449_rtl_pc = spc449_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(449*4)]   <= 1'b0;
                  active_thread[(449*4)+1] <= 1'b0;
                  active_thread[(449*4)+2] <= 1'b0;
                  active_thread[(449*4)+3] <= 1'b0;
                  spc449_inst_done         <= 0;
                  spc449_phy_pc_w          <= 0;
                end else begin
                  active_thread[(449*4)]   <= 1'b1;
                  active_thread[(449*4)+1] <= 1'b1;
                  active_thread[(449*4)+2] <= 1'b1;
                  active_thread[(449*4)+3] <= 1'b1;
                  spc449_inst_done         <= `ARIANE_CORE449.piton_pc_vld;
                  spc449_phy_pc_w          <= `ARIANE_CORE449.piton_pc;
                end
            end
    

            assign spc450_thread_id = 2'b00;
            assign spc450_rtl_pc = spc450_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(450*4)]   <= 1'b0;
                  active_thread[(450*4)+1] <= 1'b0;
                  active_thread[(450*4)+2] <= 1'b0;
                  active_thread[(450*4)+3] <= 1'b0;
                  spc450_inst_done         <= 0;
                  spc450_phy_pc_w          <= 0;
                end else begin
                  active_thread[(450*4)]   <= 1'b1;
                  active_thread[(450*4)+1] <= 1'b1;
                  active_thread[(450*4)+2] <= 1'b1;
                  active_thread[(450*4)+3] <= 1'b1;
                  spc450_inst_done         <= `ARIANE_CORE450.piton_pc_vld;
                  spc450_phy_pc_w          <= `ARIANE_CORE450.piton_pc;
                end
            end
    

            assign spc451_thread_id = 2'b00;
            assign spc451_rtl_pc = spc451_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(451*4)]   <= 1'b0;
                  active_thread[(451*4)+1] <= 1'b0;
                  active_thread[(451*4)+2] <= 1'b0;
                  active_thread[(451*4)+3] <= 1'b0;
                  spc451_inst_done         <= 0;
                  spc451_phy_pc_w          <= 0;
                end else begin
                  active_thread[(451*4)]   <= 1'b1;
                  active_thread[(451*4)+1] <= 1'b1;
                  active_thread[(451*4)+2] <= 1'b1;
                  active_thread[(451*4)+3] <= 1'b1;
                  spc451_inst_done         <= `ARIANE_CORE451.piton_pc_vld;
                  spc451_phy_pc_w          <= `ARIANE_CORE451.piton_pc;
                end
            end
    

            assign spc452_thread_id = 2'b00;
            assign spc452_rtl_pc = spc452_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(452*4)]   <= 1'b0;
                  active_thread[(452*4)+1] <= 1'b0;
                  active_thread[(452*4)+2] <= 1'b0;
                  active_thread[(452*4)+3] <= 1'b0;
                  spc452_inst_done         <= 0;
                  spc452_phy_pc_w          <= 0;
                end else begin
                  active_thread[(452*4)]   <= 1'b1;
                  active_thread[(452*4)+1] <= 1'b1;
                  active_thread[(452*4)+2] <= 1'b1;
                  active_thread[(452*4)+3] <= 1'b1;
                  spc452_inst_done         <= `ARIANE_CORE452.piton_pc_vld;
                  spc452_phy_pc_w          <= `ARIANE_CORE452.piton_pc;
                end
            end
    

            assign spc453_thread_id = 2'b00;
            assign spc453_rtl_pc = spc453_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(453*4)]   <= 1'b0;
                  active_thread[(453*4)+1] <= 1'b0;
                  active_thread[(453*4)+2] <= 1'b0;
                  active_thread[(453*4)+3] <= 1'b0;
                  spc453_inst_done         <= 0;
                  spc453_phy_pc_w          <= 0;
                end else begin
                  active_thread[(453*4)]   <= 1'b1;
                  active_thread[(453*4)+1] <= 1'b1;
                  active_thread[(453*4)+2] <= 1'b1;
                  active_thread[(453*4)+3] <= 1'b1;
                  spc453_inst_done         <= `ARIANE_CORE453.piton_pc_vld;
                  spc453_phy_pc_w          <= `ARIANE_CORE453.piton_pc;
                end
            end
    

            assign spc454_thread_id = 2'b00;
            assign spc454_rtl_pc = spc454_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(454*4)]   <= 1'b0;
                  active_thread[(454*4)+1] <= 1'b0;
                  active_thread[(454*4)+2] <= 1'b0;
                  active_thread[(454*4)+3] <= 1'b0;
                  spc454_inst_done         <= 0;
                  spc454_phy_pc_w          <= 0;
                end else begin
                  active_thread[(454*4)]   <= 1'b1;
                  active_thread[(454*4)+1] <= 1'b1;
                  active_thread[(454*4)+2] <= 1'b1;
                  active_thread[(454*4)+3] <= 1'b1;
                  spc454_inst_done         <= `ARIANE_CORE454.piton_pc_vld;
                  spc454_phy_pc_w          <= `ARIANE_CORE454.piton_pc;
                end
            end
    

            assign spc455_thread_id = 2'b00;
            assign spc455_rtl_pc = spc455_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(455*4)]   <= 1'b0;
                  active_thread[(455*4)+1] <= 1'b0;
                  active_thread[(455*4)+2] <= 1'b0;
                  active_thread[(455*4)+3] <= 1'b0;
                  spc455_inst_done         <= 0;
                  spc455_phy_pc_w          <= 0;
                end else begin
                  active_thread[(455*4)]   <= 1'b1;
                  active_thread[(455*4)+1] <= 1'b1;
                  active_thread[(455*4)+2] <= 1'b1;
                  active_thread[(455*4)+3] <= 1'b1;
                  spc455_inst_done         <= `ARIANE_CORE455.piton_pc_vld;
                  spc455_phy_pc_w          <= `ARIANE_CORE455.piton_pc;
                end
            end
    

            assign spc456_thread_id = 2'b00;
            assign spc456_rtl_pc = spc456_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(456*4)]   <= 1'b0;
                  active_thread[(456*4)+1] <= 1'b0;
                  active_thread[(456*4)+2] <= 1'b0;
                  active_thread[(456*4)+3] <= 1'b0;
                  spc456_inst_done         <= 0;
                  spc456_phy_pc_w          <= 0;
                end else begin
                  active_thread[(456*4)]   <= 1'b1;
                  active_thread[(456*4)+1] <= 1'b1;
                  active_thread[(456*4)+2] <= 1'b1;
                  active_thread[(456*4)+3] <= 1'b1;
                  spc456_inst_done         <= `ARIANE_CORE456.piton_pc_vld;
                  spc456_phy_pc_w          <= `ARIANE_CORE456.piton_pc;
                end
            end
    

            assign spc457_thread_id = 2'b00;
            assign spc457_rtl_pc = spc457_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(457*4)]   <= 1'b0;
                  active_thread[(457*4)+1] <= 1'b0;
                  active_thread[(457*4)+2] <= 1'b0;
                  active_thread[(457*4)+3] <= 1'b0;
                  spc457_inst_done         <= 0;
                  spc457_phy_pc_w          <= 0;
                end else begin
                  active_thread[(457*4)]   <= 1'b1;
                  active_thread[(457*4)+1] <= 1'b1;
                  active_thread[(457*4)+2] <= 1'b1;
                  active_thread[(457*4)+3] <= 1'b1;
                  spc457_inst_done         <= `ARIANE_CORE457.piton_pc_vld;
                  spc457_phy_pc_w          <= `ARIANE_CORE457.piton_pc;
                end
            end
    

            assign spc458_thread_id = 2'b00;
            assign spc458_rtl_pc = spc458_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(458*4)]   <= 1'b0;
                  active_thread[(458*4)+1] <= 1'b0;
                  active_thread[(458*4)+2] <= 1'b0;
                  active_thread[(458*4)+3] <= 1'b0;
                  spc458_inst_done         <= 0;
                  spc458_phy_pc_w          <= 0;
                end else begin
                  active_thread[(458*4)]   <= 1'b1;
                  active_thread[(458*4)+1] <= 1'b1;
                  active_thread[(458*4)+2] <= 1'b1;
                  active_thread[(458*4)+3] <= 1'b1;
                  spc458_inst_done         <= `ARIANE_CORE458.piton_pc_vld;
                  spc458_phy_pc_w          <= `ARIANE_CORE458.piton_pc;
                end
            end
    

            assign spc459_thread_id = 2'b00;
            assign spc459_rtl_pc = spc459_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(459*4)]   <= 1'b0;
                  active_thread[(459*4)+1] <= 1'b0;
                  active_thread[(459*4)+2] <= 1'b0;
                  active_thread[(459*4)+3] <= 1'b0;
                  spc459_inst_done         <= 0;
                  spc459_phy_pc_w          <= 0;
                end else begin
                  active_thread[(459*4)]   <= 1'b1;
                  active_thread[(459*4)+1] <= 1'b1;
                  active_thread[(459*4)+2] <= 1'b1;
                  active_thread[(459*4)+3] <= 1'b1;
                  spc459_inst_done         <= `ARIANE_CORE459.piton_pc_vld;
                  spc459_phy_pc_w          <= `ARIANE_CORE459.piton_pc;
                end
            end
    

            assign spc460_thread_id = 2'b00;
            assign spc460_rtl_pc = spc460_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(460*4)]   <= 1'b0;
                  active_thread[(460*4)+1] <= 1'b0;
                  active_thread[(460*4)+2] <= 1'b0;
                  active_thread[(460*4)+3] <= 1'b0;
                  spc460_inst_done         <= 0;
                  spc460_phy_pc_w          <= 0;
                end else begin
                  active_thread[(460*4)]   <= 1'b1;
                  active_thread[(460*4)+1] <= 1'b1;
                  active_thread[(460*4)+2] <= 1'b1;
                  active_thread[(460*4)+3] <= 1'b1;
                  spc460_inst_done         <= `ARIANE_CORE460.piton_pc_vld;
                  spc460_phy_pc_w          <= `ARIANE_CORE460.piton_pc;
                end
            end
    

            assign spc461_thread_id = 2'b00;
            assign spc461_rtl_pc = spc461_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(461*4)]   <= 1'b0;
                  active_thread[(461*4)+1] <= 1'b0;
                  active_thread[(461*4)+2] <= 1'b0;
                  active_thread[(461*4)+3] <= 1'b0;
                  spc461_inst_done         <= 0;
                  spc461_phy_pc_w          <= 0;
                end else begin
                  active_thread[(461*4)]   <= 1'b1;
                  active_thread[(461*4)+1] <= 1'b1;
                  active_thread[(461*4)+2] <= 1'b1;
                  active_thread[(461*4)+3] <= 1'b1;
                  spc461_inst_done         <= `ARIANE_CORE461.piton_pc_vld;
                  spc461_phy_pc_w          <= `ARIANE_CORE461.piton_pc;
                end
            end
    

            assign spc462_thread_id = 2'b00;
            assign spc462_rtl_pc = spc462_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(462*4)]   <= 1'b0;
                  active_thread[(462*4)+1] <= 1'b0;
                  active_thread[(462*4)+2] <= 1'b0;
                  active_thread[(462*4)+3] <= 1'b0;
                  spc462_inst_done         <= 0;
                  spc462_phy_pc_w          <= 0;
                end else begin
                  active_thread[(462*4)]   <= 1'b1;
                  active_thread[(462*4)+1] <= 1'b1;
                  active_thread[(462*4)+2] <= 1'b1;
                  active_thread[(462*4)+3] <= 1'b1;
                  spc462_inst_done         <= `ARIANE_CORE462.piton_pc_vld;
                  spc462_phy_pc_w          <= `ARIANE_CORE462.piton_pc;
                end
            end
    

            assign spc463_thread_id = 2'b00;
            assign spc463_rtl_pc = spc463_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(463*4)]   <= 1'b0;
                  active_thread[(463*4)+1] <= 1'b0;
                  active_thread[(463*4)+2] <= 1'b0;
                  active_thread[(463*4)+3] <= 1'b0;
                  spc463_inst_done         <= 0;
                  spc463_phy_pc_w          <= 0;
                end else begin
                  active_thread[(463*4)]   <= 1'b1;
                  active_thread[(463*4)+1] <= 1'b1;
                  active_thread[(463*4)+2] <= 1'b1;
                  active_thread[(463*4)+3] <= 1'b1;
                  spc463_inst_done         <= `ARIANE_CORE463.piton_pc_vld;
                  spc463_phy_pc_w          <= `ARIANE_CORE463.piton_pc;
                end
            end
    

            assign spc464_thread_id = 2'b00;
            assign spc464_rtl_pc = spc464_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(464*4)]   <= 1'b0;
                  active_thread[(464*4)+1] <= 1'b0;
                  active_thread[(464*4)+2] <= 1'b0;
                  active_thread[(464*4)+3] <= 1'b0;
                  spc464_inst_done         <= 0;
                  spc464_phy_pc_w          <= 0;
                end else begin
                  active_thread[(464*4)]   <= 1'b1;
                  active_thread[(464*4)+1] <= 1'b1;
                  active_thread[(464*4)+2] <= 1'b1;
                  active_thread[(464*4)+3] <= 1'b1;
                  spc464_inst_done         <= `ARIANE_CORE464.piton_pc_vld;
                  spc464_phy_pc_w          <= `ARIANE_CORE464.piton_pc;
                end
            end
    

            assign spc465_thread_id = 2'b00;
            assign spc465_rtl_pc = spc465_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(465*4)]   <= 1'b0;
                  active_thread[(465*4)+1] <= 1'b0;
                  active_thread[(465*4)+2] <= 1'b0;
                  active_thread[(465*4)+3] <= 1'b0;
                  spc465_inst_done         <= 0;
                  spc465_phy_pc_w          <= 0;
                end else begin
                  active_thread[(465*4)]   <= 1'b1;
                  active_thread[(465*4)+1] <= 1'b1;
                  active_thread[(465*4)+2] <= 1'b1;
                  active_thread[(465*4)+3] <= 1'b1;
                  spc465_inst_done         <= `ARIANE_CORE465.piton_pc_vld;
                  spc465_phy_pc_w          <= `ARIANE_CORE465.piton_pc;
                end
            end
    

            assign spc466_thread_id = 2'b00;
            assign spc466_rtl_pc = spc466_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(466*4)]   <= 1'b0;
                  active_thread[(466*4)+1] <= 1'b0;
                  active_thread[(466*4)+2] <= 1'b0;
                  active_thread[(466*4)+3] <= 1'b0;
                  spc466_inst_done         <= 0;
                  spc466_phy_pc_w          <= 0;
                end else begin
                  active_thread[(466*4)]   <= 1'b1;
                  active_thread[(466*4)+1] <= 1'b1;
                  active_thread[(466*4)+2] <= 1'b1;
                  active_thread[(466*4)+3] <= 1'b1;
                  spc466_inst_done         <= `ARIANE_CORE466.piton_pc_vld;
                  spc466_phy_pc_w          <= `ARIANE_CORE466.piton_pc;
                end
            end
    

            assign spc467_thread_id = 2'b00;
            assign spc467_rtl_pc = spc467_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(467*4)]   <= 1'b0;
                  active_thread[(467*4)+1] <= 1'b0;
                  active_thread[(467*4)+2] <= 1'b0;
                  active_thread[(467*4)+3] <= 1'b0;
                  spc467_inst_done         <= 0;
                  spc467_phy_pc_w          <= 0;
                end else begin
                  active_thread[(467*4)]   <= 1'b1;
                  active_thread[(467*4)+1] <= 1'b1;
                  active_thread[(467*4)+2] <= 1'b1;
                  active_thread[(467*4)+3] <= 1'b1;
                  spc467_inst_done         <= `ARIANE_CORE467.piton_pc_vld;
                  spc467_phy_pc_w          <= `ARIANE_CORE467.piton_pc;
                end
            end
    

            assign spc468_thread_id = 2'b00;
            assign spc468_rtl_pc = spc468_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(468*4)]   <= 1'b0;
                  active_thread[(468*4)+1] <= 1'b0;
                  active_thread[(468*4)+2] <= 1'b0;
                  active_thread[(468*4)+3] <= 1'b0;
                  spc468_inst_done         <= 0;
                  spc468_phy_pc_w          <= 0;
                end else begin
                  active_thread[(468*4)]   <= 1'b1;
                  active_thread[(468*4)+1] <= 1'b1;
                  active_thread[(468*4)+2] <= 1'b1;
                  active_thread[(468*4)+3] <= 1'b1;
                  spc468_inst_done         <= `ARIANE_CORE468.piton_pc_vld;
                  spc468_phy_pc_w          <= `ARIANE_CORE468.piton_pc;
                end
            end
    

            assign spc469_thread_id = 2'b00;
            assign spc469_rtl_pc = spc469_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(469*4)]   <= 1'b0;
                  active_thread[(469*4)+1] <= 1'b0;
                  active_thread[(469*4)+2] <= 1'b0;
                  active_thread[(469*4)+3] <= 1'b0;
                  spc469_inst_done         <= 0;
                  spc469_phy_pc_w          <= 0;
                end else begin
                  active_thread[(469*4)]   <= 1'b1;
                  active_thread[(469*4)+1] <= 1'b1;
                  active_thread[(469*4)+2] <= 1'b1;
                  active_thread[(469*4)+3] <= 1'b1;
                  spc469_inst_done         <= `ARIANE_CORE469.piton_pc_vld;
                  spc469_phy_pc_w          <= `ARIANE_CORE469.piton_pc;
                end
            end
    

            assign spc470_thread_id = 2'b00;
            assign spc470_rtl_pc = spc470_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(470*4)]   <= 1'b0;
                  active_thread[(470*4)+1] <= 1'b0;
                  active_thread[(470*4)+2] <= 1'b0;
                  active_thread[(470*4)+3] <= 1'b0;
                  spc470_inst_done         <= 0;
                  spc470_phy_pc_w          <= 0;
                end else begin
                  active_thread[(470*4)]   <= 1'b1;
                  active_thread[(470*4)+1] <= 1'b1;
                  active_thread[(470*4)+2] <= 1'b1;
                  active_thread[(470*4)+3] <= 1'b1;
                  spc470_inst_done         <= `ARIANE_CORE470.piton_pc_vld;
                  spc470_phy_pc_w          <= `ARIANE_CORE470.piton_pc;
                end
            end
    

            assign spc471_thread_id = 2'b00;
            assign spc471_rtl_pc = spc471_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(471*4)]   <= 1'b0;
                  active_thread[(471*4)+1] <= 1'b0;
                  active_thread[(471*4)+2] <= 1'b0;
                  active_thread[(471*4)+3] <= 1'b0;
                  spc471_inst_done         <= 0;
                  spc471_phy_pc_w          <= 0;
                end else begin
                  active_thread[(471*4)]   <= 1'b1;
                  active_thread[(471*4)+1] <= 1'b1;
                  active_thread[(471*4)+2] <= 1'b1;
                  active_thread[(471*4)+3] <= 1'b1;
                  spc471_inst_done         <= `ARIANE_CORE471.piton_pc_vld;
                  spc471_phy_pc_w          <= `ARIANE_CORE471.piton_pc;
                end
            end
    

            assign spc472_thread_id = 2'b00;
            assign spc472_rtl_pc = spc472_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(472*4)]   <= 1'b0;
                  active_thread[(472*4)+1] <= 1'b0;
                  active_thread[(472*4)+2] <= 1'b0;
                  active_thread[(472*4)+3] <= 1'b0;
                  spc472_inst_done         <= 0;
                  spc472_phy_pc_w          <= 0;
                end else begin
                  active_thread[(472*4)]   <= 1'b1;
                  active_thread[(472*4)+1] <= 1'b1;
                  active_thread[(472*4)+2] <= 1'b1;
                  active_thread[(472*4)+3] <= 1'b1;
                  spc472_inst_done         <= `ARIANE_CORE472.piton_pc_vld;
                  spc472_phy_pc_w          <= `ARIANE_CORE472.piton_pc;
                end
            end
    

            assign spc473_thread_id = 2'b00;
            assign spc473_rtl_pc = spc473_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(473*4)]   <= 1'b0;
                  active_thread[(473*4)+1] <= 1'b0;
                  active_thread[(473*4)+2] <= 1'b0;
                  active_thread[(473*4)+3] <= 1'b0;
                  spc473_inst_done         <= 0;
                  spc473_phy_pc_w          <= 0;
                end else begin
                  active_thread[(473*4)]   <= 1'b1;
                  active_thread[(473*4)+1] <= 1'b1;
                  active_thread[(473*4)+2] <= 1'b1;
                  active_thread[(473*4)+3] <= 1'b1;
                  spc473_inst_done         <= `ARIANE_CORE473.piton_pc_vld;
                  spc473_phy_pc_w          <= `ARIANE_CORE473.piton_pc;
                end
            end
    

            assign spc474_thread_id = 2'b00;
            assign spc474_rtl_pc = spc474_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(474*4)]   <= 1'b0;
                  active_thread[(474*4)+1] <= 1'b0;
                  active_thread[(474*4)+2] <= 1'b0;
                  active_thread[(474*4)+3] <= 1'b0;
                  spc474_inst_done         <= 0;
                  spc474_phy_pc_w          <= 0;
                end else begin
                  active_thread[(474*4)]   <= 1'b1;
                  active_thread[(474*4)+1] <= 1'b1;
                  active_thread[(474*4)+2] <= 1'b1;
                  active_thread[(474*4)+3] <= 1'b1;
                  spc474_inst_done         <= `ARIANE_CORE474.piton_pc_vld;
                  spc474_phy_pc_w          <= `ARIANE_CORE474.piton_pc;
                end
            end
    

            assign spc475_thread_id = 2'b00;
            assign spc475_rtl_pc = spc475_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(475*4)]   <= 1'b0;
                  active_thread[(475*4)+1] <= 1'b0;
                  active_thread[(475*4)+2] <= 1'b0;
                  active_thread[(475*4)+3] <= 1'b0;
                  spc475_inst_done         <= 0;
                  spc475_phy_pc_w          <= 0;
                end else begin
                  active_thread[(475*4)]   <= 1'b1;
                  active_thread[(475*4)+1] <= 1'b1;
                  active_thread[(475*4)+2] <= 1'b1;
                  active_thread[(475*4)+3] <= 1'b1;
                  spc475_inst_done         <= `ARIANE_CORE475.piton_pc_vld;
                  spc475_phy_pc_w          <= `ARIANE_CORE475.piton_pc;
                end
            end
    

            assign spc476_thread_id = 2'b00;
            assign spc476_rtl_pc = spc476_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(476*4)]   <= 1'b0;
                  active_thread[(476*4)+1] <= 1'b0;
                  active_thread[(476*4)+2] <= 1'b0;
                  active_thread[(476*4)+3] <= 1'b0;
                  spc476_inst_done         <= 0;
                  spc476_phy_pc_w          <= 0;
                end else begin
                  active_thread[(476*4)]   <= 1'b1;
                  active_thread[(476*4)+1] <= 1'b1;
                  active_thread[(476*4)+2] <= 1'b1;
                  active_thread[(476*4)+3] <= 1'b1;
                  spc476_inst_done         <= `ARIANE_CORE476.piton_pc_vld;
                  spc476_phy_pc_w          <= `ARIANE_CORE476.piton_pc;
                end
            end
    

            assign spc477_thread_id = 2'b00;
            assign spc477_rtl_pc = spc477_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(477*4)]   <= 1'b0;
                  active_thread[(477*4)+1] <= 1'b0;
                  active_thread[(477*4)+2] <= 1'b0;
                  active_thread[(477*4)+3] <= 1'b0;
                  spc477_inst_done         <= 0;
                  spc477_phy_pc_w          <= 0;
                end else begin
                  active_thread[(477*4)]   <= 1'b1;
                  active_thread[(477*4)+1] <= 1'b1;
                  active_thread[(477*4)+2] <= 1'b1;
                  active_thread[(477*4)+3] <= 1'b1;
                  spc477_inst_done         <= `ARIANE_CORE477.piton_pc_vld;
                  spc477_phy_pc_w          <= `ARIANE_CORE477.piton_pc;
                end
            end
    

            assign spc478_thread_id = 2'b00;
            assign spc478_rtl_pc = spc478_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(478*4)]   <= 1'b0;
                  active_thread[(478*4)+1] <= 1'b0;
                  active_thread[(478*4)+2] <= 1'b0;
                  active_thread[(478*4)+3] <= 1'b0;
                  spc478_inst_done         <= 0;
                  spc478_phy_pc_w          <= 0;
                end else begin
                  active_thread[(478*4)]   <= 1'b1;
                  active_thread[(478*4)+1] <= 1'b1;
                  active_thread[(478*4)+2] <= 1'b1;
                  active_thread[(478*4)+3] <= 1'b1;
                  spc478_inst_done         <= `ARIANE_CORE478.piton_pc_vld;
                  spc478_phy_pc_w          <= `ARIANE_CORE478.piton_pc;
                end
            end
    

            assign spc479_thread_id = 2'b00;
            assign spc479_rtl_pc = spc479_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(479*4)]   <= 1'b0;
                  active_thread[(479*4)+1] <= 1'b0;
                  active_thread[(479*4)+2] <= 1'b0;
                  active_thread[(479*4)+3] <= 1'b0;
                  spc479_inst_done         <= 0;
                  spc479_phy_pc_w          <= 0;
                end else begin
                  active_thread[(479*4)]   <= 1'b1;
                  active_thread[(479*4)+1] <= 1'b1;
                  active_thread[(479*4)+2] <= 1'b1;
                  active_thread[(479*4)+3] <= 1'b1;
                  spc479_inst_done         <= `ARIANE_CORE479.piton_pc_vld;
                  spc479_phy_pc_w          <= `ARIANE_CORE479.piton_pc;
                end
            end
    

            assign spc480_thread_id = 2'b00;
            assign spc480_rtl_pc = spc480_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(480*4)]   <= 1'b0;
                  active_thread[(480*4)+1] <= 1'b0;
                  active_thread[(480*4)+2] <= 1'b0;
                  active_thread[(480*4)+3] <= 1'b0;
                  spc480_inst_done         <= 0;
                  spc480_phy_pc_w          <= 0;
                end else begin
                  active_thread[(480*4)]   <= 1'b1;
                  active_thread[(480*4)+1] <= 1'b1;
                  active_thread[(480*4)+2] <= 1'b1;
                  active_thread[(480*4)+3] <= 1'b1;
                  spc480_inst_done         <= `ARIANE_CORE480.piton_pc_vld;
                  spc480_phy_pc_w          <= `ARIANE_CORE480.piton_pc;
                end
            end
    

            assign spc481_thread_id = 2'b00;
            assign spc481_rtl_pc = spc481_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(481*4)]   <= 1'b0;
                  active_thread[(481*4)+1] <= 1'b0;
                  active_thread[(481*4)+2] <= 1'b0;
                  active_thread[(481*4)+3] <= 1'b0;
                  spc481_inst_done         <= 0;
                  spc481_phy_pc_w          <= 0;
                end else begin
                  active_thread[(481*4)]   <= 1'b1;
                  active_thread[(481*4)+1] <= 1'b1;
                  active_thread[(481*4)+2] <= 1'b1;
                  active_thread[(481*4)+3] <= 1'b1;
                  spc481_inst_done         <= `ARIANE_CORE481.piton_pc_vld;
                  spc481_phy_pc_w          <= `ARIANE_CORE481.piton_pc;
                end
            end
    

            assign spc482_thread_id = 2'b00;
            assign spc482_rtl_pc = spc482_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(482*4)]   <= 1'b0;
                  active_thread[(482*4)+1] <= 1'b0;
                  active_thread[(482*4)+2] <= 1'b0;
                  active_thread[(482*4)+3] <= 1'b0;
                  spc482_inst_done         <= 0;
                  spc482_phy_pc_w          <= 0;
                end else begin
                  active_thread[(482*4)]   <= 1'b1;
                  active_thread[(482*4)+1] <= 1'b1;
                  active_thread[(482*4)+2] <= 1'b1;
                  active_thread[(482*4)+3] <= 1'b1;
                  spc482_inst_done         <= `ARIANE_CORE482.piton_pc_vld;
                  spc482_phy_pc_w          <= `ARIANE_CORE482.piton_pc;
                end
            end
    

            assign spc483_thread_id = 2'b00;
            assign spc483_rtl_pc = spc483_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(483*4)]   <= 1'b0;
                  active_thread[(483*4)+1] <= 1'b0;
                  active_thread[(483*4)+2] <= 1'b0;
                  active_thread[(483*4)+3] <= 1'b0;
                  spc483_inst_done         <= 0;
                  spc483_phy_pc_w          <= 0;
                end else begin
                  active_thread[(483*4)]   <= 1'b1;
                  active_thread[(483*4)+1] <= 1'b1;
                  active_thread[(483*4)+2] <= 1'b1;
                  active_thread[(483*4)+3] <= 1'b1;
                  spc483_inst_done         <= `ARIANE_CORE483.piton_pc_vld;
                  spc483_phy_pc_w          <= `ARIANE_CORE483.piton_pc;
                end
            end
    

            assign spc484_thread_id = 2'b00;
            assign spc484_rtl_pc = spc484_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(484*4)]   <= 1'b0;
                  active_thread[(484*4)+1] <= 1'b0;
                  active_thread[(484*4)+2] <= 1'b0;
                  active_thread[(484*4)+3] <= 1'b0;
                  spc484_inst_done         <= 0;
                  spc484_phy_pc_w          <= 0;
                end else begin
                  active_thread[(484*4)]   <= 1'b1;
                  active_thread[(484*4)+1] <= 1'b1;
                  active_thread[(484*4)+2] <= 1'b1;
                  active_thread[(484*4)+3] <= 1'b1;
                  spc484_inst_done         <= `ARIANE_CORE484.piton_pc_vld;
                  spc484_phy_pc_w          <= `ARIANE_CORE484.piton_pc;
                end
            end
    

            assign spc485_thread_id = 2'b00;
            assign spc485_rtl_pc = spc485_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(485*4)]   <= 1'b0;
                  active_thread[(485*4)+1] <= 1'b0;
                  active_thread[(485*4)+2] <= 1'b0;
                  active_thread[(485*4)+3] <= 1'b0;
                  spc485_inst_done         <= 0;
                  spc485_phy_pc_w          <= 0;
                end else begin
                  active_thread[(485*4)]   <= 1'b1;
                  active_thread[(485*4)+1] <= 1'b1;
                  active_thread[(485*4)+2] <= 1'b1;
                  active_thread[(485*4)+3] <= 1'b1;
                  spc485_inst_done         <= `ARIANE_CORE485.piton_pc_vld;
                  spc485_phy_pc_w          <= `ARIANE_CORE485.piton_pc;
                end
            end
    

            assign spc486_thread_id = 2'b00;
            assign spc486_rtl_pc = spc486_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(486*4)]   <= 1'b0;
                  active_thread[(486*4)+1] <= 1'b0;
                  active_thread[(486*4)+2] <= 1'b0;
                  active_thread[(486*4)+3] <= 1'b0;
                  spc486_inst_done         <= 0;
                  spc486_phy_pc_w          <= 0;
                end else begin
                  active_thread[(486*4)]   <= 1'b1;
                  active_thread[(486*4)+1] <= 1'b1;
                  active_thread[(486*4)+2] <= 1'b1;
                  active_thread[(486*4)+3] <= 1'b1;
                  spc486_inst_done         <= `ARIANE_CORE486.piton_pc_vld;
                  spc486_phy_pc_w          <= `ARIANE_CORE486.piton_pc;
                end
            end
    

            assign spc487_thread_id = 2'b00;
            assign spc487_rtl_pc = spc487_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(487*4)]   <= 1'b0;
                  active_thread[(487*4)+1] <= 1'b0;
                  active_thread[(487*4)+2] <= 1'b0;
                  active_thread[(487*4)+3] <= 1'b0;
                  spc487_inst_done         <= 0;
                  spc487_phy_pc_w          <= 0;
                end else begin
                  active_thread[(487*4)]   <= 1'b1;
                  active_thread[(487*4)+1] <= 1'b1;
                  active_thread[(487*4)+2] <= 1'b1;
                  active_thread[(487*4)+3] <= 1'b1;
                  spc487_inst_done         <= `ARIANE_CORE487.piton_pc_vld;
                  spc487_phy_pc_w          <= `ARIANE_CORE487.piton_pc;
                end
            end
    

            assign spc488_thread_id = 2'b00;
            assign spc488_rtl_pc = spc488_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(488*4)]   <= 1'b0;
                  active_thread[(488*4)+1] <= 1'b0;
                  active_thread[(488*4)+2] <= 1'b0;
                  active_thread[(488*4)+3] <= 1'b0;
                  spc488_inst_done         <= 0;
                  spc488_phy_pc_w          <= 0;
                end else begin
                  active_thread[(488*4)]   <= 1'b1;
                  active_thread[(488*4)+1] <= 1'b1;
                  active_thread[(488*4)+2] <= 1'b1;
                  active_thread[(488*4)+3] <= 1'b1;
                  spc488_inst_done         <= `ARIANE_CORE488.piton_pc_vld;
                  spc488_phy_pc_w          <= `ARIANE_CORE488.piton_pc;
                end
            end
    

            assign spc489_thread_id = 2'b00;
            assign spc489_rtl_pc = spc489_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(489*4)]   <= 1'b0;
                  active_thread[(489*4)+1] <= 1'b0;
                  active_thread[(489*4)+2] <= 1'b0;
                  active_thread[(489*4)+3] <= 1'b0;
                  spc489_inst_done         <= 0;
                  spc489_phy_pc_w          <= 0;
                end else begin
                  active_thread[(489*4)]   <= 1'b1;
                  active_thread[(489*4)+1] <= 1'b1;
                  active_thread[(489*4)+2] <= 1'b1;
                  active_thread[(489*4)+3] <= 1'b1;
                  spc489_inst_done         <= `ARIANE_CORE489.piton_pc_vld;
                  spc489_phy_pc_w          <= `ARIANE_CORE489.piton_pc;
                end
            end
    

            assign spc490_thread_id = 2'b00;
            assign spc490_rtl_pc = spc490_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(490*4)]   <= 1'b0;
                  active_thread[(490*4)+1] <= 1'b0;
                  active_thread[(490*4)+2] <= 1'b0;
                  active_thread[(490*4)+3] <= 1'b0;
                  spc490_inst_done         <= 0;
                  spc490_phy_pc_w          <= 0;
                end else begin
                  active_thread[(490*4)]   <= 1'b1;
                  active_thread[(490*4)+1] <= 1'b1;
                  active_thread[(490*4)+2] <= 1'b1;
                  active_thread[(490*4)+3] <= 1'b1;
                  spc490_inst_done         <= `ARIANE_CORE490.piton_pc_vld;
                  spc490_phy_pc_w          <= `ARIANE_CORE490.piton_pc;
                end
            end
    

            assign spc491_thread_id = 2'b00;
            assign spc491_rtl_pc = spc491_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(491*4)]   <= 1'b0;
                  active_thread[(491*4)+1] <= 1'b0;
                  active_thread[(491*4)+2] <= 1'b0;
                  active_thread[(491*4)+3] <= 1'b0;
                  spc491_inst_done         <= 0;
                  spc491_phy_pc_w          <= 0;
                end else begin
                  active_thread[(491*4)]   <= 1'b1;
                  active_thread[(491*4)+1] <= 1'b1;
                  active_thread[(491*4)+2] <= 1'b1;
                  active_thread[(491*4)+3] <= 1'b1;
                  spc491_inst_done         <= `ARIANE_CORE491.piton_pc_vld;
                  spc491_phy_pc_w          <= `ARIANE_CORE491.piton_pc;
                end
            end
    

            assign spc492_thread_id = 2'b00;
            assign spc492_rtl_pc = spc492_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(492*4)]   <= 1'b0;
                  active_thread[(492*4)+1] <= 1'b0;
                  active_thread[(492*4)+2] <= 1'b0;
                  active_thread[(492*4)+3] <= 1'b0;
                  spc492_inst_done         <= 0;
                  spc492_phy_pc_w          <= 0;
                end else begin
                  active_thread[(492*4)]   <= 1'b1;
                  active_thread[(492*4)+1] <= 1'b1;
                  active_thread[(492*4)+2] <= 1'b1;
                  active_thread[(492*4)+3] <= 1'b1;
                  spc492_inst_done         <= `ARIANE_CORE492.piton_pc_vld;
                  spc492_phy_pc_w          <= `ARIANE_CORE492.piton_pc;
                end
            end
    

            assign spc493_thread_id = 2'b00;
            assign spc493_rtl_pc = spc493_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(493*4)]   <= 1'b0;
                  active_thread[(493*4)+1] <= 1'b0;
                  active_thread[(493*4)+2] <= 1'b0;
                  active_thread[(493*4)+3] <= 1'b0;
                  spc493_inst_done         <= 0;
                  spc493_phy_pc_w          <= 0;
                end else begin
                  active_thread[(493*4)]   <= 1'b1;
                  active_thread[(493*4)+1] <= 1'b1;
                  active_thread[(493*4)+2] <= 1'b1;
                  active_thread[(493*4)+3] <= 1'b1;
                  spc493_inst_done         <= `ARIANE_CORE493.piton_pc_vld;
                  spc493_phy_pc_w          <= `ARIANE_CORE493.piton_pc;
                end
            end
    

            assign spc494_thread_id = 2'b00;
            assign spc494_rtl_pc = spc494_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(494*4)]   <= 1'b0;
                  active_thread[(494*4)+1] <= 1'b0;
                  active_thread[(494*4)+2] <= 1'b0;
                  active_thread[(494*4)+3] <= 1'b0;
                  spc494_inst_done         <= 0;
                  spc494_phy_pc_w          <= 0;
                end else begin
                  active_thread[(494*4)]   <= 1'b1;
                  active_thread[(494*4)+1] <= 1'b1;
                  active_thread[(494*4)+2] <= 1'b1;
                  active_thread[(494*4)+3] <= 1'b1;
                  spc494_inst_done         <= `ARIANE_CORE494.piton_pc_vld;
                  spc494_phy_pc_w          <= `ARIANE_CORE494.piton_pc;
                end
            end
    

            assign spc495_thread_id = 2'b00;
            assign spc495_rtl_pc = spc495_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(495*4)]   <= 1'b0;
                  active_thread[(495*4)+1] <= 1'b0;
                  active_thread[(495*4)+2] <= 1'b0;
                  active_thread[(495*4)+3] <= 1'b0;
                  spc495_inst_done         <= 0;
                  spc495_phy_pc_w          <= 0;
                end else begin
                  active_thread[(495*4)]   <= 1'b1;
                  active_thread[(495*4)+1] <= 1'b1;
                  active_thread[(495*4)+2] <= 1'b1;
                  active_thread[(495*4)+3] <= 1'b1;
                  spc495_inst_done         <= `ARIANE_CORE495.piton_pc_vld;
                  spc495_phy_pc_w          <= `ARIANE_CORE495.piton_pc;
                end
            end
    

            assign spc496_thread_id = 2'b00;
            assign spc496_rtl_pc = spc496_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(496*4)]   <= 1'b0;
                  active_thread[(496*4)+1] <= 1'b0;
                  active_thread[(496*4)+2] <= 1'b0;
                  active_thread[(496*4)+3] <= 1'b0;
                  spc496_inst_done         <= 0;
                  spc496_phy_pc_w          <= 0;
                end else begin
                  active_thread[(496*4)]   <= 1'b1;
                  active_thread[(496*4)+1] <= 1'b1;
                  active_thread[(496*4)+2] <= 1'b1;
                  active_thread[(496*4)+3] <= 1'b1;
                  spc496_inst_done         <= `ARIANE_CORE496.piton_pc_vld;
                  spc496_phy_pc_w          <= `ARIANE_CORE496.piton_pc;
                end
            end
    

            assign spc497_thread_id = 2'b00;
            assign spc497_rtl_pc = spc497_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(497*4)]   <= 1'b0;
                  active_thread[(497*4)+1] <= 1'b0;
                  active_thread[(497*4)+2] <= 1'b0;
                  active_thread[(497*4)+3] <= 1'b0;
                  spc497_inst_done         <= 0;
                  spc497_phy_pc_w          <= 0;
                end else begin
                  active_thread[(497*4)]   <= 1'b1;
                  active_thread[(497*4)+1] <= 1'b1;
                  active_thread[(497*4)+2] <= 1'b1;
                  active_thread[(497*4)+3] <= 1'b1;
                  spc497_inst_done         <= `ARIANE_CORE497.piton_pc_vld;
                  spc497_phy_pc_w          <= `ARIANE_CORE497.piton_pc;
                end
            end
    

            assign spc498_thread_id = 2'b00;
            assign spc498_rtl_pc = spc498_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(498*4)]   <= 1'b0;
                  active_thread[(498*4)+1] <= 1'b0;
                  active_thread[(498*4)+2] <= 1'b0;
                  active_thread[(498*4)+3] <= 1'b0;
                  spc498_inst_done         <= 0;
                  spc498_phy_pc_w          <= 0;
                end else begin
                  active_thread[(498*4)]   <= 1'b1;
                  active_thread[(498*4)+1] <= 1'b1;
                  active_thread[(498*4)+2] <= 1'b1;
                  active_thread[(498*4)+3] <= 1'b1;
                  spc498_inst_done         <= `ARIANE_CORE498.piton_pc_vld;
                  spc498_phy_pc_w          <= `ARIANE_CORE498.piton_pc;
                end
            end
    

            assign spc499_thread_id = 2'b00;
            assign spc499_rtl_pc = spc499_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(499*4)]   <= 1'b0;
                  active_thread[(499*4)+1] <= 1'b0;
                  active_thread[(499*4)+2] <= 1'b0;
                  active_thread[(499*4)+3] <= 1'b0;
                  spc499_inst_done         <= 0;
                  spc499_phy_pc_w          <= 0;
                end else begin
                  active_thread[(499*4)]   <= 1'b1;
                  active_thread[(499*4)+1] <= 1'b1;
                  active_thread[(499*4)+2] <= 1'b1;
                  active_thread[(499*4)+3] <= 1'b1;
                  spc499_inst_done         <= `ARIANE_CORE499.piton_pc_vld;
                  spc499_phy_pc_w          <= `ARIANE_CORE499.piton_pc;
                end
            end
    

            assign spc500_thread_id = 2'b00;
            assign spc500_rtl_pc = spc500_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(500*4)]   <= 1'b0;
                  active_thread[(500*4)+1] <= 1'b0;
                  active_thread[(500*4)+2] <= 1'b0;
                  active_thread[(500*4)+3] <= 1'b0;
                  spc500_inst_done         <= 0;
                  spc500_phy_pc_w          <= 0;
                end else begin
                  active_thread[(500*4)]   <= 1'b1;
                  active_thread[(500*4)+1] <= 1'b1;
                  active_thread[(500*4)+2] <= 1'b1;
                  active_thread[(500*4)+3] <= 1'b1;
                  spc500_inst_done         <= `ARIANE_CORE500.piton_pc_vld;
                  spc500_phy_pc_w          <= `ARIANE_CORE500.piton_pc;
                end
            end
    

            assign spc501_thread_id = 2'b00;
            assign spc501_rtl_pc = spc501_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(501*4)]   <= 1'b0;
                  active_thread[(501*4)+1] <= 1'b0;
                  active_thread[(501*4)+2] <= 1'b0;
                  active_thread[(501*4)+3] <= 1'b0;
                  spc501_inst_done         <= 0;
                  spc501_phy_pc_w          <= 0;
                end else begin
                  active_thread[(501*4)]   <= 1'b1;
                  active_thread[(501*4)+1] <= 1'b1;
                  active_thread[(501*4)+2] <= 1'b1;
                  active_thread[(501*4)+3] <= 1'b1;
                  spc501_inst_done         <= `ARIANE_CORE501.piton_pc_vld;
                  spc501_phy_pc_w          <= `ARIANE_CORE501.piton_pc;
                end
            end
    

            assign spc502_thread_id = 2'b00;
            assign spc502_rtl_pc = spc502_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(502*4)]   <= 1'b0;
                  active_thread[(502*4)+1] <= 1'b0;
                  active_thread[(502*4)+2] <= 1'b0;
                  active_thread[(502*4)+3] <= 1'b0;
                  spc502_inst_done         <= 0;
                  spc502_phy_pc_w          <= 0;
                end else begin
                  active_thread[(502*4)]   <= 1'b1;
                  active_thread[(502*4)+1] <= 1'b1;
                  active_thread[(502*4)+2] <= 1'b1;
                  active_thread[(502*4)+3] <= 1'b1;
                  spc502_inst_done         <= `ARIANE_CORE502.piton_pc_vld;
                  spc502_phy_pc_w          <= `ARIANE_CORE502.piton_pc;
                end
            end
    

            assign spc503_thread_id = 2'b00;
            assign spc503_rtl_pc = spc503_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(503*4)]   <= 1'b0;
                  active_thread[(503*4)+1] <= 1'b0;
                  active_thread[(503*4)+2] <= 1'b0;
                  active_thread[(503*4)+3] <= 1'b0;
                  spc503_inst_done         <= 0;
                  spc503_phy_pc_w          <= 0;
                end else begin
                  active_thread[(503*4)]   <= 1'b1;
                  active_thread[(503*4)+1] <= 1'b1;
                  active_thread[(503*4)+2] <= 1'b1;
                  active_thread[(503*4)+3] <= 1'b1;
                  spc503_inst_done         <= `ARIANE_CORE503.piton_pc_vld;
                  spc503_phy_pc_w          <= `ARIANE_CORE503.piton_pc;
                end
            end
    

            assign spc504_thread_id = 2'b00;
            assign spc504_rtl_pc = spc504_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(504*4)]   <= 1'b0;
                  active_thread[(504*4)+1] <= 1'b0;
                  active_thread[(504*4)+2] <= 1'b0;
                  active_thread[(504*4)+3] <= 1'b0;
                  spc504_inst_done         <= 0;
                  spc504_phy_pc_w          <= 0;
                end else begin
                  active_thread[(504*4)]   <= 1'b1;
                  active_thread[(504*4)+1] <= 1'b1;
                  active_thread[(504*4)+2] <= 1'b1;
                  active_thread[(504*4)+3] <= 1'b1;
                  spc504_inst_done         <= `ARIANE_CORE504.piton_pc_vld;
                  spc504_phy_pc_w          <= `ARIANE_CORE504.piton_pc;
                end
            end
    

            assign spc505_thread_id = 2'b00;
            assign spc505_rtl_pc = spc505_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(505*4)]   <= 1'b0;
                  active_thread[(505*4)+1] <= 1'b0;
                  active_thread[(505*4)+2] <= 1'b0;
                  active_thread[(505*4)+3] <= 1'b0;
                  spc505_inst_done         <= 0;
                  spc505_phy_pc_w          <= 0;
                end else begin
                  active_thread[(505*4)]   <= 1'b1;
                  active_thread[(505*4)+1] <= 1'b1;
                  active_thread[(505*4)+2] <= 1'b1;
                  active_thread[(505*4)+3] <= 1'b1;
                  spc505_inst_done         <= `ARIANE_CORE505.piton_pc_vld;
                  spc505_phy_pc_w          <= `ARIANE_CORE505.piton_pc;
                end
            end
    

            assign spc506_thread_id = 2'b00;
            assign spc506_rtl_pc = spc506_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(506*4)]   <= 1'b0;
                  active_thread[(506*4)+1] <= 1'b0;
                  active_thread[(506*4)+2] <= 1'b0;
                  active_thread[(506*4)+3] <= 1'b0;
                  spc506_inst_done         <= 0;
                  spc506_phy_pc_w          <= 0;
                end else begin
                  active_thread[(506*4)]   <= 1'b1;
                  active_thread[(506*4)+1] <= 1'b1;
                  active_thread[(506*4)+2] <= 1'b1;
                  active_thread[(506*4)+3] <= 1'b1;
                  spc506_inst_done         <= `ARIANE_CORE506.piton_pc_vld;
                  spc506_phy_pc_w          <= `ARIANE_CORE506.piton_pc;
                end
            end
    

            assign spc507_thread_id = 2'b00;
            assign spc507_rtl_pc = spc507_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(507*4)]   <= 1'b0;
                  active_thread[(507*4)+1] <= 1'b0;
                  active_thread[(507*4)+2] <= 1'b0;
                  active_thread[(507*4)+3] <= 1'b0;
                  spc507_inst_done         <= 0;
                  spc507_phy_pc_w          <= 0;
                end else begin
                  active_thread[(507*4)]   <= 1'b1;
                  active_thread[(507*4)+1] <= 1'b1;
                  active_thread[(507*4)+2] <= 1'b1;
                  active_thread[(507*4)+3] <= 1'b1;
                  spc507_inst_done         <= `ARIANE_CORE507.piton_pc_vld;
                  spc507_phy_pc_w          <= `ARIANE_CORE507.piton_pc;
                end
            end
    

            assign spc508_thread_id = 2'b00;
            assign spc508_rtl_pc = spc508_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(508*4)]   <= 1'b0;
                  active_thread[(508*4)+1] <= 1'b0;
                  active_thread[(508*4)+2] <= 1'b0;
                  active_thread[(508*4)+3] <= 1'b0;
                  spc508_inst_done         <= 0;
                  spc508_phy_pc_w          <= 0;
                end else begin
                  active_thread[(508*4)]   <= 1'b1;
                  active_thread[(508*4)+1] <= 1'b1;
                  active_thread[(508*4)+2] <= 1'b1;
                  active_thread[(508*4)+3] <= 1'b1;
                  spc508_inst_done         <= `ARIANE_CORE508.piton_pc_vld;
                  spc508_phy_pc_w          <= `ARIANE_CORE508.piton_pc;
                end
            end
    

            assign spc509_thread_id = 2'b00;
            assign spc509_rtl_pc = spc509_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(509*4)]   <= 1'b0;
                  active_thread[(509*4)+1] <= 1'b0;
                  active_thread[(509*4)+2] <= 1'b0;
                  active_thread[(509*4)+3] <= 1'b0;
                  spc509_inst_done         <= 0;
                  spc509_phy_pc_w          <= 0;
                end else begin
                  active_thread[(509*4)]   <= 1'b1;
                  active_thread[(509*4)+1] <= 1'b1;
                  active_thread[(509*4)+2] <= 1'b1;
                  active_thread[(509*4)+3] <= 1'b1;
                  spc509_inst_done         <= `ARIANE_CORE509.piton_pc_vld;
                  spc509_phy_pc_w          <= `ARIANE_CORE509.piton_pc;
                end
            end
    

            assign spc510_thread_id = 2'b00;
            assign spc510_rtl_pc = spc510_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(510*4)]   <= 1'b0;
                  active_thread[(510*4)+1] <= 1'b0;
                  active_thread[(510*4)+2] <= 1'b0;
                  active_thread[(510*4)+3] <= 1'b0;
                  spc510_inst_done         <= 0;
                  spc510_phy_pc_w          <= 0;
                end else begin
                  active_thread[(510*4)]   <= 1'b1;
                  active_thread[(510*4)+1] <= 1'b1;
                  active_thread[(510*4)+2] <= 1'b1;
                  active_thread[(510*4)+3] <= 1'b1;
                  spc510_inst_done         <= `ARIANE_CORE510.piton_pc_vld;
                  spc510_phy_pc_w          <= `ARIANE_CORE510.piton_pc;
                end
            end
    

            assign spc511_thread_id = 2'b00;
            assign spc511_rtl_pc = spc511_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(511*4)]   <= 1'b0;
                  active_thread[(511*4)+1] <= 1'b0;
                  active_thread[(511*4)+2] <= 1'b0;
                  active_thread[(511*4)+3] <= 1'b0;
                  spc511_inst_done         <= 0;
                  spc511_phy_pc_w          <= 0;
                end else begin
                  active_thread[(511*4)]   <= 1'b1;
                  active_thread[(511*4)+1] <= 1'b1;
                  active_thread[(511*4)+2] <= 1'b1;
                  active_thread[(511*4)+3] <= 1'b1;
                  spc511_inst_done         <= `ARIANE_CORE511.piton_pc_vld;
                  spc511_phy_pc_w          <= `ARIANE_CORE511.piton_pc;
                end
            end
    

            assign spc512_thread_id = 2'b00;
            assign spc512_rtl_pc = spc512_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(512*4)]   <= 1'b0;
                  active_thread[(512*4)+1] <= 1'b0;
                  active_thread[(512*4)+2] <= 1'b0;
                  active_thread[(512*4)+3] <= 1'b0;
                  spc512_inst_done         <= 0;
                  spc512_phy_pc_w          <= 0;
                end else begin
                  active_thread[(512*4)]   <= 1'b1;
                  active_thread[(512*4)+1] <= 1'b1;
                  active_thread[(512*4)+2] <= 1'b1;
                  active_thread[(512*4)+3] <= 1'b1;
                  spc512_inst_done         <= `ARIANE_CORE512.piton_pc_vld;
                  spc512_phy_pc_w          <= `ARIANE_CORE512.piton_pc;
                end
            end
    

            assign spc513_thread_id = 2'b00;
            assign spc513_rtl_pc = spc513_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(513*4)]   <= 1'b0;
                  active_thread[(513*4)+1] <= 1'b0;
                  active_thread[(513*4)+2] <= 1'b0;
                  active_thread[(513*4)+3] <= 1'b0;
                  spc513_inst_done         <= 0;
                  spc513_phy_pc_w          <= 0;
                end else begin
                  active_thread[(513*4)]   <= 1'b1;
                  active_thread[(513*4)+1] <= 1'b1;
                  active_thread[(513*4)+2] <= 1'b1;
                  active_thread[(513*4)+3] <= 1'b1;
                  spc513_inst_done         <= `ARIANE_CORE513.piton_pc_vld;
                  spc513_phy_pc_w          <= `ARIANE_CORE513.piton_pc;
                end
            end
    

            assign spc514_thread_id = 2'b00;
            assign spc514_rtl_pc = spc514_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(514*4)]   <= 1'b0;
                  active_thread[(514*4)+1] <= 1'b0;
                  active_thread[(514*4)+2] <= 1'b0;
                  active_thread[(514*4)+3] <= 1'b0;
                  spc514_inst_done         <= 0;
                  spc514_phy_pc_w          <= 0;
                end else begin
                  active_thread[(514*4)]   <= 1'b1;
                  active_thread[(514*4)+1] <= 1'b1;
                  active_thread[(514*4)+2] <= 1'b1;
                  active_thread[(514*4)+3] <= 1'b1;
                  spc514_inst_done         <= `ARIANE_CORE514.piton_pc_vld;
                  spc514_phy_pc_w          <= `ARIANE_CORE514.piton_pc;
                end
            end
    

            assign spc515_thread_id = 2'b00;
            assign spc515_rtl_pc = spc515_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(515*4)]   <= 1'b0;
                  active_thread[(515*4)+1] <= 1'b0;
                  active_thread[(515*4)+2] <= 1'b0;
                  active_thread[(515*4)+3] <= 1'b0;
                  spc515_inst_done         <= 0;
                  spc515_phy_pc_w          <= 0;
                end else begin
                  active_thread[(515*4)]   <= 1'b1;
                  active_thread[(515*4)+1] <= 1'b1;
                  active_thread[(515*4)+2] <= 1'b1;
                  active_thread[(515*4)+3] <= 1'b1;
                  spc515_inst_done         <= `ARIANE_CORE515.piton_pc_vld;
                  spc515_phy_pc_w          <= `ARIANE_CORE515.piton_pc;
                end
            end
    

            assign spc516_thread_id = 2'b00;
            assign spc516_rtl_pc = spc516_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(516*4)]   <= 1'b0;
                  active_thread[(516*4)+1] <= 1'b0;
                  active_thread[(516*4)+2] <= 1'b0;
                  active_thread[(516*4)+3] <= 1'b0;
                  spc516_inst_done         <= 0;
                  spc516_phy_pc_w          <= 0;
                end else begin
                  active_thread[(516*4)]   <= 1'b1;
                  active_thread[(516*4)+1] <= 1'b1;
                  active_thread[(516*4)+2] <= 1'b1;
                  active_thread[(516*4)+3] <= 1'b1;
                  spc516_inst_done         <= `ARIANE_CORE516.piton_pc_vld;
                  spc516_phy_pc_w          <= `ARIANE_CORE516.piton_pc;
                end
            end
    

            assign spc517_thread_id = 2'b00;
            assign spc517_rtl_pc = spc517_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(517*4)]   <= 1'b0;
                  active_thread[(517*4)+1] <= 1'b0;
                  active_thread[(517*4)+2] <= 1'b0;
                  active_thread[(517*4)+3] <= 1'b0;
                  spc517_inst_done         <= 0;
                  spc517_phy_pc_w          <= 0;
                end else begin
                  active_thread[(517*4)]   <= 1'b1;
                  active_thread[(517*4)+1] <= 1'b1;
                  active_thread[(517*4)+2] <= 1'b1;
                  active_thread[(517*4)+3] <= 1'b1;
                  spc517_inst_done         <= `ARIANE_CORE517.piton_pc_vld;
                  spc517_phy_pc_w          <= `ARIANE_CORE517.piton_pc;
                end
            end
    

            assign spc518_thread_id = 2'b00;
            assign spc518_rtl_pc = spc518_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(518*4)]   <= 1'b0;
                  active_thread[(518*4)+1] <= 1'b0;
                  active_thread[(518*4)+2] <= 1'b0;
                  active_thread[(518*4)+3] <= 1'b0;
                  spc518_inst_done         <= 0;
                  spc518_phy_pc_w          <= 0;
                end else begin
                  active_thread[(518*4)]   <= 1'b1;
                  active_thread[(518*4)+1] <= 1'b1;
                  active_thread[(518*4)+2] <= 1'b1;
                  active_thread[(518*4)+3] <= 1'b1;
                  spc518_inst_done         <= `ARIANE_CORE518.piton_pc_vld;
                  spc518_phy_pc_w          <= `ARIANE_CORE518.piton_pc;
                end
            end
    

            assign spc519_thread_id = 2'b00;
            assign spc519_rtl_pc = spc519_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(519*4)]   <= 1'b0;
                  active_thread[(519*4)+1] <= 1'b0;
                  active_thread[(519*4)+2] <= 1'b0;
                  active_thread[(519*4)+3] <= 1'b0;
                  spc519_inst_done         <= 0;
                  spc519_phy_pc_w          <= 0;
                end else begin
                  active_thread[(519*4)]   <= 1'b1;
                  active_thread[(519*4)+1] <= 1'b1;
                  active_thread[(519*4)+2] <= 1'b1;
                  active_thread[(519*4)+3] <= 1'b1;
                  spc519_inst_done         <= `ARIANE_CORE519.piton_pc_vld;
                  spc519_phy_pc_w          <= `ARIANE_CORE519.piton_pc;
                end
            end
    

            assign spc520_thread_id = 2'b00;
            assign spc520_rtl_pc = spc520_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(520*4)]   <= 1'b0;
                  active_thread[(520*4)+1] <= 1'b0;
                  active_thread[(520*4)+2] <= 1'b0;
                  active_thread[(520*4)+3] <= 1'b0;
                  spc520_inst_done         <= 0;
                  spc520_phy_pc_w          <= 0;
                end else begin
                  active_thread[(520*4)]   <= 1'b1;
                  active_thread[(520*4)+1] <= 1'b1;
                  active_thread[(520*4)+2] <= 1'b1;
                  active_thread[(520*4)+3] <= 1'b1;
                  spc520_inst_done         <= `ARIANE_CORE520.piton_pc_vld;
                  spc520_phy_pc_w          <= `ARIANE_CORE520.piton_pc;
                end
            end
    

            assign spc521_thread_id = 2'b00;
            assign spc521_rtl_pc = spc521_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(521*4)]   <= 1'b0;
                  active_thread[(521*4)+1] <= 1'b0;
                  active_thread[(521*4)+2] <= 1'b0;
                  active_thread[(521*4)+3] <= 1'b0;
                  spc521_inst_done         <= 0;
                  spc521_phy_pc_w          <= 0;
                end else begin
                  active_thread[(521*4)]   <= 1'b1;
                  active_thread[(521*4)+1] <= 1'b1;
                  active_thread[(521*4)+2] <= 1'b1;
                  active_thread[(521*4)+3] <= 1'b1;
                  spc521_inst_done         <= `ARIANE_CORE521.piton_pc_vld;
                  spc521_phy_pc_w          <= `ARIANE_CORE521.piton_pc;
                end
            end
    

            assign spc522_thread_id = 2'b00;
            assign spc522_rtl_pc = spc522_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(522*4)]   <= 1'b0;
                  active_thread[(522*4)+1] <= 1'b0;
                  active_thread[(522*4)+2] <= 1'b0;
                  active_thread[(522*4)+3] <= 1'b0;
                  spc522_inst_done         <= 0;
                  spc522_phy_pc_w          <= 0;
                end else begin
                  active_thread[(522*4)]   <= 1'b1;
                  active_thread[(522*4)+1] <= 1'b1;
                  active_thread[(522*4)+2] <= 1'b1;
                  active_thread[(522*4)+3] <= 1'b1;
                  spc522_inst_done         <= `ARIANE_CORE522.piton_pc_vld;
                  spc522_phy_pc_w          <= `ARIANE_CORE522.piton_pc;
                end
            end
    

            assign spc523_thread_id = 2'b00;
            assign spc523_rtl_pc = spc523_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(523*4)]   <= 1'b0;
                  active_thread[(523*4)+1] <= 1'b0;
                  active_thread[(523*4)+2] <= 1'b0;
                  active_thread[(523*4)+3] <= 1'b0;
                  spc523_inst_done         <= 0;
                  spc523_phy_pc_w          <= 0;
                end else begin
                  active_thread[(523*4)]   <= 1'b1;
                  active_thread[(523*4)+1] <= 1'b1;
                  active_thread[(523*4)+2] <= 1'b1;
                  active_thread[(523*4)+3] <= 1'b1;
                  spc523_inst_done         <= `ARIANE_CORE523.piton_pc_vld;
                  spc523_phy_pc_w          <= `ARIANE_CORE523.piton_pc;
                end
            end
    

            assign spc524_thread_id = 2'b00;
            assign spc524_rtl_pc = spc524_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(524*4)]   <= 1'b0;
                  active_thread[(524*4)+1] <= 1'b0;
                  active_thread[(524*4)+2] <= 1'b0;
                  active_thread[(524*4)+3] <= 1'b0;
                  spc524_inst_done         <= 0;
                  spc524_phy_pc_w          <= 0;
                end else begin
                  active_thread[(524*4)]   <= 1'b1;
                  active_thread[(524*4)+1] <= 1'b1;
                  active_thread[(524*4)+2] <= 1'b1;
                  active_thread[(524*4)+3] <= 1'b1;
                  spc524_inst_done         <= `ARIANE_CORE524.piton_pc_vld;
                  spc524_phy_pc_w          <= `ARIANE_CORE524.piton_pc;
                end
            end
    

            assign spc525_thread_id = 2'b00;
            assign spc525_rtl_pc = spc525_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(525*4)]   <= 1'b0;
                  active_thread[(525*4)+1] <= 1'b0;
                  active_thread[(525*4)+2] <= 1'b0;
                  active_thread[(525*4)+3] <= 1'b0;
                  spc525_inst_done         <= 0;
                  spc525_phy_pc_w          <= 0;
                end else begin
                  active_thread[(525*4)]   <= 1'b1;
                  active_thread[(525*4)+1] <= 1'b1;
                  active_thread[(525*4)+2] <= 1'b1;
                  active_thread[(525*4)+3] <= 1'b1;
                  spc525_inst_done         <= `ARIANE_CORE525.piton_pc_vld;
                  spc525_phy_pc_w          <= `ARIANE_CORE525.piton_pc;
                end
            end
    

            assign spc526_thread_id = 2'b00;
            assign spc526_rtl_pc = spc526_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(526*4)]   <= 1'b0;
                  active_thread[(526*4)+1] <= 1'b0;
                  active_thread[(526*4)+2] <= 1'b0;
                  active_thread[(526*4)+3] <= 1'b0;
                  spc526_inst_done         <= 0;
                  spc526_phy_pc_w          <= 0;
                end else begin
                  active_thread[(526*4)]   <= 1'b1;
                  active_thread[(526*4)+1] <= 1'b1;
                  active_thread[(526*4)+2] <= 1'b1;
                  active_thread[(526*4)+3] <= 1'b1;
                  spc526_inst_done         <= `ARIANE_CORE526.piton_pc_vld;
                  spc526_phy_pc_w          <= `ARIANE_CORE526.piton_pc;
                end
            end
    

            assign spc527_thread_id = 2'b00;
            assign spc527_rtl_pc = spc527_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(527*4)]   <= 1'b0;
                  active_thread[(527*4)+1] <= 1'b0;
                  active_thread[(527*4)+2] <= 1'b0;
                  active_thread[(527*4)+3] <= 1'b0;
                  spc527_inst_done         <= 0;
                  spc527_phy_pc_w          <= 0;
                end else begin
                  active_thread[(527*4)]   <= 1'b1;
                  active_thread[(527*4)+1] <= 1'b1;
                  active_thread[(527*4)+2] <= 1'b1;
                  active_thread[(527*4)+3] <= 1'b1;
                  spc527_inst_done         <= `ARIANE_CORE527.piton_pc_vld;
                  spc527_phy_pc_w          <= `ARIANE_CORE527.piton_pc;
                end
            end
    

            assign spc528_thread_id = 2'b00;
            assign spc528_rtl_pc = spc528_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(528*4)]   <= 1'b0;
                  active_thread[(528*4)+1] <= 1'b0;
                  active_thread[(528*4)+2] <= 1'b0;
                  active_thread[(528*4)+3] <= 1'b0;
                  spc528_inst_done         <= 0;
                  spc528_phy_pc_w          <= 0;
                end else begin
                  active_thread[(528*4)]   <= 1'b1;
                  active_thread[(528*4)+1] <= 1'b1;
                  active_thread[(528*4)+2] <= 1'b1;
                  active_thread[(528*4)+3] <= 1'b1;
                  spc528_inst_done         <= `ARIANE_CORE528.piton_pc_vld;
                  spc528_phy_pc_w          <= `ARIANE_CORE528.piton_pc;
                end
            end
    

            assign spc529_thread_id = 2'b00;
            assign spc529_rtl_pc = spc529_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(529*4)]   <= 1'b0;
                  active_thread[(529*4)+1] <= 1'b0;
                  active_thread[(529*4)+2] <= 1'b0;
                  active_thread[(529*4)+3] <= 1'b0;
                  spc529_inst_done         <= 0;
                  spc529_phy_pc_w          <= 0;
                end else begin
                  active_thread[(529*4)]   <= 1'b1;
                  active_thread[(529*4)+1] <= 1'b1;
                  active_thread[(529*4)+2] <= 1'b1;
                  active_thread[(529*4)+3] <= 1'b1;
                  spc529_inst_done         <= `ARIANE_CORE529.piton_pc_vld;
                  spc529_phy_pc_w          <= `ARIANE_CORE529.piton_pc;
                end
            end
    

            assign spc530_thread_id = 2'b00;
            assign spc530_rtl_pc = spc530_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(530*4)]   <= 1'b0;
                  active_thread[(530*4)+1] <= 1'b0;
                  active_thread[(530*4)+2] <= 1'b0;
                  active_thread[(530*4)+3] <= 1'b0;
                  spc530_inst_done         <= 0;
                  spc530_phy_pc_w          <= 0;
                end else begin
                  active_thread[(530*4)]   <= 1'b1;
                  active_thread[(530*4)+1] <= 1'b1;
                  active_thread[(530*4)+2] <= 1'b1;
                  active_thread[(530*4)+3] <= 1'b1;
                  spc530_inst_done         <= `ARIANE_CORE530.piton_pc_vld;
                  spc530_phy_pc_w          <= `ARIANE_CORE530.piton_pc;
                end
            end
    

            assign spc531_thread_id = 2'b00;
            assign spc531_rtl_pc = spc531_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(531*4)]   <= 1'b0;
                  active_thread[(531*4)+1] <= 1'b0;
                  active_thread[(531*4)+2] <= 1'b0;
                  active_thread[(531*4)+3] <= 1'b0;
                  spc531_inst_done         <= 0;
                  spc531_phy_pc_w          <= 0;
                end else begin
                  active_thread[(531*4)]   <= 1'b1;
                  active_thread[(531*4)+1] <= 1'b1;
                  active_thread[(531*4)+2] <= 1'b1;
                  active_thread[(531*4)+3] <= 1'b1;
                  spc531_inst_done         <= `ARIANE_CORE531.piton_pc_vld;
                  spc531_phy_pc_w          <= `ARIANE_CORE531.piton_pc;
                end
            end
    

            assign spc532_thread_id = 2'b00;
            assign spc532_rtl_pc = spc532_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(532*4)]   <= 1'b0;
                  active_thread[(532*4)+1] <= 1'b0;
                  active_thread[(532*4)+2] <= 1'b0;
                  active_thread[(532*4)+3] <= 1'b0;
                  spc532_inst_done         <= 0;
                  spc532_phy_pc_w          <= 0;
                end else begin
                  active_thread[(532*4)]   <= 1'b1;
                  active_thread[(532*4)+1] <= 1'b1;
                  active_thread[(532*4)+2] <= 1'b1;
                  active_thread[(532*4)+3] <= 1'b1;
                  spc532_inst_done         <= `ARIANE_CORE532.piton_pc_vld;
                  spc532_phy_pc_w          <= `ARIANE_CORE532.piton_pc;
                end
            end
    

            assign spc533_thread_id = 2'b00;
            assign spc533_rtl_pc = spc533_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(533*4)]   <= 1'b0;
                  active_thread[(533*4)+1] <= 1'b0;
                  active_thread[(533*4)+2] <= 1'b0;
                  active_thread[(533*4)+3] <= 1'b0;
                  spc533_inst_done         <= 0;
                  spc533_phy_pc_w          <= 0;
                end else begin
                  active_thread[(533*4)]   <= 1'b1;
                  active_thread[(533*4)+1] <= 1'b1;
                  active_thread[(533*4)+2] <= 1'b1;
                  active_thread[(533*4)+3] <= 1'b1;
                  spc533_inst_done         <= `ARIANE_CORE533.piton_pc_vld;
                  spc533_phy_pc_w          <= `ARIANE_CORE533.piton_pc;
                end
            end
    

            assign spc534_thread_id = 2'b00;
            assign spc534_rtl_pc = spc534_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(534*4)]   <= 1'b0;
                  active_thread[(534*4)+1] <= 1'b0;
                  active_thread[(534*4)+2] <= 1'b0;
                  active_thread[(534*4)+3] <= 1'b0;
                  spc534_inst_done         <= 0;
                  spc534_phy_pc_w          <= 0;
                end else begin
                  active_thread[(534*4)]   <= 1'b1;
                  active_thread[(534*4)+1] <= 1'b1;
                  active_thread[(534*4)+2] <= 1'b1;
                  active_thread[(534*4)+3] <= 1'b1;
                  spc534_inst_done         <= `ARIANE_CORE534.piton_pc_vld;
                  spc534_phy_pc_w          <= `ARIANE_CORE534.piton_pc;
                end
            end
    

            assign spc535_thread_id = 2'b00;
            assign spc535_rtl_pc = spc535_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(535*4)]   <= 1'b0;
                  active_thread[(535*4)+1] <= 1'b0;
                  active_thread[(535*4)+2] <= 1'b0;
                  active_thread[(535*4)+3] <= 1'b0;
                  spc535_inst_done         <= 0;
                  spc535_phy_pc_w          <= 0;
                end else begin
                  active_thread[(535*4)]   <= 1'b1;
                  active_thread[(535*4)+1] <= 1'b1;
                  active_thread[(535*4)+2] <= 1'b1;
                  active_thread[(535*4)+3] <= 1'b1;
                  spc535_inst_done         <= `ARIANE_CORE535.piton_pc_vld;
                  spc535_phy_pc_w          <= `ARIANE_CORE535.piton_pc;
                end
            end
    

            assign spc536_thread_id = 2'b00;
            assign spc536_rtl_pc = spc536_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(536*4)]   <= 1'b0;
                  active_thread[(536*4)+1] <= 1'b0;
                  active_thread[(536*4)+2] <= 1'b0;
                  active_thread[(536*4)+3] <= 1'b0;
                  spc536_inst_done         <= 0;
                  spc536_phy_pc_w          <= 0;
                end else begin
                  active_thread[(536*4)]   <= 1'b1;
                  active_thread[(536*4)+1] <= 1'b1;
                  active_thread[(536*4)+2] <= 1'b1;
                  active_thread[(536*4)+3] <= 1'b1;
                  spc536_inst_done         <= `ARIANE_CORE536.piton_pc_vld;
                  spc536_phy_pc_w          <= `ARIANE_CORE536.piton_pc;
                end
            end
    

            assign spc537_thread_id = 2'b00;
            assign spc537_rtl_pc = spc537_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(537*4)]   <= 1'b0;
                  active_thread[(537*4)+1] <= 1'b0;
                  active_thread[(537*4)+2] <= 1'b0;
                  active_thread[(537*4)+3] <= 1'b0;
                  spc537_inst_done         <= 0;
                  spc537_phy_pc_w          <= 0;
                end else begin
                  active_thread[(537*4)]   <= 1'b1;
                  active_thread[(537*4)+1] <= 1'b1;
                  active_thread[(537*4)+2] <= 1'b1;
                  active_thread[(537*4)+3] <= 1'b1;
                  spc537_inst_done         <= `ARIANE_CORE537.piton_pc_vld;
                  spc537_phy_pc_w          <= `ARIANE_CORE537.piton_pc;
                end
            end
    

            assign spc538_thread_id = 2'b00;
            assign spc538_rtl_pc = spc538_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(538*4)]   <= 1'b0;
                  active_thread[(538*4)+1] <= 1'b0;
                  active_thread[(538*4)+2] <= 1'b0;
                  active_thread[(538*4)+3] <= 1'b0;
                  spc538_inst_done         <= 0;
                  spc538_phy_pc_w          <= 0;
                end else begin
                  active_thread[(538*4)]   <= 1'b1;
                  active_thread[(538*4)+1] <= 1'b1;
                  active_thread[(538*4)+2] <= 1'b1;
                  active_thread[(538*4)+3] <= 1'b1;
                  spc538_inst_done         <= `ARIANE_CORE538.piton_pc_vld;
                  spc538_phy_pc_w          <= `ARIANE_CORE538.piton_pc;
                end
            end
    

            assign spc539_thread_id = 2'b00;
            assign spc539_rtl_pc = spc539_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(539*4)]   <= 1'b0;
                  active_thread[(539*4)+1] <= 1'b0;
                  active_thread[(539*4)+2] <= 1'b0;
                  active_thread[(539*4)+3] <= 1'b0;
                  spc539_inst_done         <= 0;
                  spc539_phy_pc_w          <= 0;
                end else begin
                  active_thread[(539*4)]   <= 1'b1;
                  active_thread[(539*4)+1] <= 1'b1;
                  active_thread[(539*4)+2] <= 1'b1;
                  active_thread[(539*4)+3] <= 1'b1;
                  spc539_inst_done         <= `ARIANE_CORE539.piton_pc_vld;
                  spc539_phy_pc_w          <= `ARIANE_CORE539.piton_pc;
                end
            end
    

            assign spc540_thread_id = 2'b00;
            assign spc540_rtl_pc = spc540_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(540*4)]   <= 1'b0;
                  active_thread[(540*4)+1] <= 1'b0;
                  active_thread[(540*4)+2] <= 1'b0;
                  active_thread[(540*4)+3] <= 1'b0;
                  spc540_inst_done         <= 0;
                  spc540_phy_pc_w          <= 0;
                end else begin
                  active_thread[(540*4)]   <= 1'b1;
                  active_thread[(540*4)+1] <= 1'b1;
                  active_thread[(540*4)+2] <= 1'b1;
                  active_thread[(540*4)+3] <= 1'b1;
                  spc540_inst_done         <= `ARIANE_CORE540.piton_pc_vld;
                  spc540_phy_pc_w          <= `ARIANE_CORE540.piton_pc;
                end
            end
    

            assign spc541_thread_id = 2'b00;
            assign spc541_rtl_pc = spc541_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(541*4)]   <= 1'b0;
                  active_thread[(541*4)+1] <= 1'b0;
                  active_thread[(541*4)+2] <= 1'b0;
                  active_thread[(541*4)+3] <= 1'b0;
                  spc541_inst_done         <= 0;
                  spc541_phy_pc_w          <= 0;
                end else begin
                  active_thread[(541*4)]   <= 1'b1;
                  active_thread[(541*4)+1] <= 1'b1;
                  active_thread[(541*4)+2] <= 1'b1;
                  active_thread[(541*4)+3] <= 1'b1;
                  spc541_inst_done         <= `ARIANE_CORE541.piton_pc_vld;
                  spc541_phy_pc_w          <= `ARIANE_CORE541.piton_pc;
                end
            end
    

            assign spc542_thread_id = 2'b00;
            assign spc542_rtl_pc = spc542_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(542*4)]   <= 1'b0;
                  active_thread[(542*4)+1] <= 1'b0;
                  active_thread[(542*4)+2] <= 1'b0;
                  active_thread[(542*4)+3] <= 1'b0;
                  spc542_inst_done         <= 0;
                  spc542_phy_pc_w          <= 0;
                end else begin
                  active_thread[(542*4)]   <= 1'b1;
                  active_thread[(542*4)+1] <= 1'b1;
                  active_thread[(542*4)+2] <= 1'b1;
                  active_thread[(542*4)+3] <= 1'b1;
                  spc542_inst_done         <= `ARIANE_CORE542.piton_pc_vld;
                  spc542_phy_pc_w          <= `ARIANE_CORE542.piton_pc;
                end
            end
    

            assign spc543_thread_id = 2'b00;
            assign spc543_rtl_pc = spc543_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(543*4)]   <= 1'b0;
                  active_thread[(543*4)+1] <= 1'b0;
                  active_thread[(543*4)+2] <= 1'b0;
                  active_thread[(543*4)+3] <= 1'b0;
                  spc543_inst_done         <= 0;
                  spc543_phy_pc_w          <= 0;
                end else begin
                  active_thread[(543*4)]   <= 1'b1;
                  active_thread[(543*4)+1] <= 1'b1;
                  active_thread[(543*4)+2] <= 1'b1;
                  active_thread[(543*4)+3] <= 1'b1;
                  spc543_inst_done         <= `ARIANE_CORE543.piton_pc_vld;
                  spc543_phy_pc_w          <= `ARIANE_CORE543.piton_pc;
                end
            end
    

            assign spc544_thread_id = 2'b00;
            assign spc544_rtl_pc = spc544_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(544*4)]   <= 1'b0;
                  active_thread[(544*4)+1] <= 1'b0;
                  active_thread[(544*4)+2] <= 1'b0;
                  active_thread[(544*4)+3] <= 1'b0;
                  spc544_inst_done         <= 0;
                  spc544_phy_pc_w          <= 0;
                end else begin
                  active_thread[(544*4)]   <= 1'b1;
                  active_thread[(544*4)+1] <= 1'b1;
                  active_thread[(544*4)+2] <= 1'b1;
                  active_thread[(544*4)+3] <= 1'b1;
                  spc544_inst_done         <= `ARIANE_CORE544.piton_pc_vld;
                  spc544_phy_pc_w          <= `ARIANE_CORE544.piton_pc;
                end
            end
    

            assign spc545_thread_id = 2'b00;
            assign spc545_rtl_pc = spc545_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(545*4)]   <= 1'b0;
                  active_thread[(545*4)+1] <= 1'b0;
                  active_thread[(545*4)+2] <= 1'b0;
                  active_thread[(545*4)+3] <= 1'b0;
                  spc545_inst_done         <= 0;
                  spc545_phy_pc_w          <= 0;
                end else begin
                  active_thread[(545*4)]   <= 1'b1;
                  active_thread[(545*4)+1] <= 1'b1;
                  active_thread[(545*4)+2] <= 1'b1;
                  active_thread[(545*4)+3] <= 1'b1;
                  spc545_inst_done         <= `ARIANE_CORE545.piton_pc_vld;
                  spc545_phy_pc_w          <= `ARIANE_CORE545.piton_pc;
                end
            end
    

            assign spc546_thread_id = 2'b00;
            assign spc546_rtl_pc = spc546_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(546*4)]   <= 1'b0;
                  active_thread[(546*4)+1] <= 1'b0;
                  active_thread[(546*4)+2] <= 1'b0;
                  active_thread[(546*4)+3] <= 1'b0;
                  spc546_inst_done         <= 0;
                  spc546_phy_pc_w          <= 0;
                end else begin
                  active_thread[(546*4)]   <= 1'b1;
                  active_thread[(546*4)+1] <= 1'b1;
                  active_thread[(546*4)+2] <= 1'b1;
                  active_thread[(546*4)+3] <= 1'b1;
                  spc546_inst_done         <= `ARIANE_CORE546.piton_pc_vld;
                  spc546_phy_pc_w          <= `ARIANE_CORE546.piton_pc;
                end
            end
    

            assign spc547_thread_id = 2'b00;
            assign spc547_rtl_pc = spc547_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(547*4)]   <= 1'b0;
                  active_thread[(547*4)+1] <= 1'b0;
                  active_thread[(547*4)+2] <= 1'b0;
                  active_thread[(547*4)+3] <= 1'b0;
                  spc547_inst_done         <= 0;
                  spc547_phy_pc_w          <= 0;
                end else begin
                  active_thread[(547*4)]   <= 1'b1;
                  active_thread[(547*4)+1] <= 1'b1;
                  active_thread[(547*4)+2] <= 1'b1;
                  active_thread[(547*4)+3] <= 1'b1;
                  spc547_inst_done         <= `ARIANE_CORE547.piton_pc_vld;
                  spc547_phy_pc_w          <= `ARIANE_CORE547.piton_pc;
                end
            end
    

            assign spc548_thread_id = 2'b00;
            assign spc548_rtl_pc = spc548_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(548*4)]   <= 1'b0;
                  active_thread[(548*4)+1] <= 1'b0;
                  active_thread[(548*4)+2] <= 1'b0;
                  active_thread[(548*4)+3] <= 1'b0;
                  spc548_inst_done         <= 0;
                  spc548_phy_pc_w          <= 0;
                end else begin
                  active_thread[(548*4)]   <= 1'b1;
                  active_thread[(548*4)+1] <= 1'b1;
                  active_thread[(548*4)+2] <= 1'b1;
                  active_thread[(548*4)+3] <= 1'b1;
                  spc548_inst_done         <= `ARIANE_CORE548.piton_pc_vld;
                  spc548_phy_pc_w          <= `ARIANE_CORE548.piton_pc;
                end
            end
    

            assign spc549_thread_id = 2'b00;
            assign spc549_rtl_pc = spc549_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(549*4)]   <= 1'b0;
                  active_thread[(549*4)+1] <= 1'b0;
                  active_thread[(549*4)+2] <= 1'b0;
                  active_thread[(549*4)+3] <= 1'b0;
                  spc549_inst_done         <= 0;
                  spc549_phy_pc_w          <= 0;
                end else begin
                  active_thread[(549*4)]   <= 1'b1;
                  active_thread[(549*4)+1] <= 1'b1;
                  active_thread[(549*4)+2] <= 1'b1;
                  active_thread[(549*4)+3] <= 1'b1;
                  spc549_inst_done         <= `ARIANE_CORE549.piton_pc_vld;
                  spc549_phy_pc_w          <= `ARIANE_CORE549.piton_pc;
                end
            end
    

            assign spc550_thread_id = 2'b00;
            assign spc550_rtl_pc = spc550_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(550*4)]   <= 1'b0;
                  active_thread[(550*4)+1] <= 1'b0;
                  active_thread[(550*4)+2] <= 1'b0;
                  active_thread[(550*4)+3] <= 1'b0;
                  spc550_inst_done         <= 0;
                  spc550_phy_pc_w          <= 0;
                end else begin
                  active_thread[(550*4)]   <= 1'b1;
                  active_thread[(550*4)+1] <= 1'b1;
                  active_thread[(550*4)+2] <= 1'b1;
                  active_thread[(550*4)+3] <= 1'b1;
                  spc550_inst_done         <= `ARIANE_CORE550.piton_pc_vld;
                  spc550_phy_pc_w          <= `ARIANE_CORE550.piton_pc;
                end
            end
    

            assign spc551_thread_id = 2'b00;
            assign spc551_rtl_pc = spc551_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(551*4)]   <= 1'b0;
                  active_thread[(551*4)+1] <= 1'b0;
                  active_thread[(551*4)+2] <= 1'b0;
                  active_thread[(551*4)+3] <= 1'b0;
                  spc551_inst_done         <= 0;
                  spc551_phy_pc_w          <= 0;
                end else begin
                  active_thread[(551*4)]   <= 1'b1;
                  active_thread[(551*4)+1] <= 1'b1;
                  active_thread[(551*4)+2] <= 1'b1;
                  active_thread[(551*4)+3] <= 1'b1;
                  spc551_inst_done         <= `ARIANE_CORE551.piton_pc_vld;
                  spc551_phy_pc_w          <= `ARIANE_CORE551.piton_pc;
                end
            end
    

            assign spc552_thread_id = 2'b00;
            assign spc552_rtl_pc = spc552_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(552*4)]   <= 1'b0;
                  active_thread[(552*4)+1] <= 1'b0;
                  active_thread[(552*4)+2] <= 1'b0;
                  active_thread[(552*4)+3] <= 1'b0;
                  spc552_inst_done         <= 0;
                  spc552_phy_pc_w          <= 0;
                end else begin
                  active_thread[(552*4)]   <= 1'b1;
                  active_thread[(552*4)+1] <= 1'b1;
                  active_thread[(552*4)+2] <= 1'b1;
                  active_thread[(552*4)+3] <= 1'b1;
                  spc552_inst_done         <= `ARIANE_CORE552.piton_pc_vld;
                  spc552_phy_pc_w          <= `ARIANE_CORE552.piton_pc;
                end
            end
    

            assign spc553_thread_id = 2'b00;
            assign spc553_rtl_pc = spc553_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(553*4)]   <= 1'b0;
                  active_thread[(553*4)+1] <= 1'b0;
                  active_thread[(553*4)+2] <= 1'b0;
                  active_thread[(553*4)+3] <= 1'b0;
                  spc553_inst_done         <= 0;
                  spc553_phy_pc_w          <= 0;
                end else begin
                  active_thread[(553*4)]   <= 1'b1;
                  active_thread[(553*4)+1] <= 1'b1;
                  active_thread[(553*4)+2] <= 1'b1;
                  active_thread[(553*4)+3] <= 1'b1;
                  spc553_inst_done         <= `ARIANE_CORE553.piton_pc_vld;
                  spc553_phy_pc_w          <= `ARIANE_CORE553.piton_pc;
                end
            end
    

            assign spc554_thread_id = 2'b00;
            assign spc554_rtl_pc = spc554_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(554*4)]   <= 1'b0;
                  active_thread[(554*4)+1] <= 1'b0;
                  active_thread[(554*4)+2] <= 1'b0;
                  active_thread[(554*4)+3] <= 1'b0;
                  spc554_inst_done         <= 0;
                  spc554_phy_pc_w          <= 0;
                end else begin
                  active_thread[(554*4)]   <= 1'b1;
                  active_thread[(554*4)+1] <= 1'b1;
                  active_thread[(554*4)+2] <= 1'b1;
                  active_thread[(554*4)+3] <= 1'b1;
                  spc554_inst_done         <= `ARIANE_CORE554.piton_pc_vld;
                  spc554_phy_pc_w          <= `ARIANE_CORE554.piton_pc;
                end
            end
    

            assign spc555_thread_id = 2'b00;
            assign spc555_rtl_pc = spc555_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(555*4)]   <= 1'b0;
                  active_thread[(555*4)+1] <= 1'b0;
                  active_thread[(555*4)+2] <= 1'b0;
                  active_thread[(555*4)+3] <= 1'b0;
                  spc555_inst_done         <= 0;
                  spc555_phy_pc_w          <= 0;
                end else begin
                  active_thread[(555*4)]   <= 1'b1;
                  active_thread[(555*4)+1] <= 1'b1;
                  active_thread[(555*4)+2] <= 1'b1;
                  active_thread[(555*4)+3] <= 1'b1;
                  spc555_inst_done         <= `ARIANE_CORE555.piton_pc_vld;
                  spc555_phy_pc_w          <= `ARIANE_CORE555.piton_pc;
                end
            end
    

            assign spc556_thread_id = 2'b00;
            assign spc556_rtl_pc = spc556_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(556*4)]   <= 1'b0;
                  active_thread[(556*4)+1] <= 1'b0;
                  active_thread[(556*4)+2] <= 1'b0;
                  active_thread[(556*4)+3] <= 1'b0;
                  spc556_inst_done         <= 0;
                  spc556_phy_pc_w          <= 0;
                end else begin
                  active_thread[(556*4)]   <= 1'b1;
                  active_thread[(556*4)+1] <= 1'b1;
                  active_thread[(556*4)+2] <= 1'b1;
                  active_thread[(556*4)+3] <= 1'b1;
                  spc556_inst_done         <= `ARIANE_CORE556.piton_pc_vld;
                  spc556_phy_pc_w          <= `ARIANE_CORE556.piton_pc;
                end
            end
    

            assign spc557_thread_id = 2'b00;
            assign spc557_rtl_pc = spc557_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(557*4)]   <= 1'b0;
                  active_thread[(557*4)+1] <= 1'b0;
                  active_thread[(557*4)+2] <= 1'b0;
                  active_thread[(557*4)+3] <= 1'b0;
                  spc557_inst_done         <= 0;
                  spc557_phy_pc_w          <= 0;
                end else begin
                  active_thread[(557*4)]   <= 1'b1;
                  active_thread[(557*4)+1] <= 1'b1;
                  active_thread[(557*4)+2] <= 1'b1;
                  active_thread[(557*4)+3] <= 1'b1;
                  spc557_inst_done         <= `ARIANE_CORE557.piton_pc_vld;
                  spc557_phy_pc_w          <= `ARIANE_CORE557.piton_pc;
                end
            end
    

            assign spc558_thread_id = 2'b00;
            assign spc558_rtl_pc = spc558_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(558*4)]   <= 1'b0;
                  active_thread[(558*4)+1] <= 1'b0;
                  active_thread[(558*4)+2] <= 1'b0;
                  active_thread[(558*4)+3] <= 1'b0;
                  spc558_inst_done         <= 0;
                  spc558_phy_pc_w          <= 0;
                end else begin
                  active_thread[(558*4)]   <= 1'b1;
                  active_thread[(558*4)+1] <= 1'b1;
                  active_thread[(558*4)+2] <= 1'b1;
                  active_thread[(558*4)+3] <= 1'b1;
                  spc558_inst_done         <= `ARIANE_CORE558.piton_pc_vld;
                  spc558_phy_pc_w          <= `ARIANE_CORE558.piton_pc;
                end
            end
    

            assign spc559_thread_id = 2'b00;
            assign spc559_rtl_pc = spc559_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(559*4)]   <= 1'b0;
                  active_thread[(559*4)+1] <= 1'b0;
                  active_thread[(559*4)+2] <= 1'b0;
                  active_thread[(559*4)+3] <= 1'b0;
                  spc559_inst_done         <= 0;
                  spc559_phy_pc_w          <= 0;
                end else begin
                  active_thread[(559*4)]   <= 1'b1;
                  active_thread[(559*4)+1] <= 1'b1;
                  active_thread[(559*4)+2] <= 1'b1;
                  active_thread[(559*4)+3] <= 1'b1;
                  spc559_inst_done         <= `ARIANE_CORE559.piton_pc_vld;
                  spc559_phy_pc_w          <= `ARIANE_CORE559.piton_pc;
                end
            end
    

            assign spc560_thread_id = 2'b00;
            assign spc560_rtl_pc = spc560_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(560*4)]   <= 1'b0;
                  active_thread[(560*4)+1] <= 1'b0;
                  active_thread[(560*4)+2] <= 1'b0;
                  active_thread[(560*4)+3] <= 1'b0;
                  spc560_inst_done         <= 0;
                  spc560_phy_pc_w          <= 0;
                end else begin
                  active_thread[(560*4)]   <= 1'b1;
                  active_thread[(560*4)+1] <= 1'b1;
                  active_thread[(560*4)+2] <= 1'b1;
                  active_thread[(560*4)+3] <= 1'b1;
                  spc560_inst_done         <= `ARIANE_CORE560.piton_pc_vld;
                  spc560_phy_pc_w          <= `ARIANE_CORE560.piton_pc;
                end
            end
    

            assign spc561_thread_id = 2'b00;
            assign spc561_rtl_pc = spc561_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(561*4)]   <= 1'b0;
                  active_thread[(561*4)+1] <= 1'b0;
                  active_thread[(561*4)+2] <= 1'b0;
                  active_thread[(561*4)+3] <= 1'b0;
                  spc561_inst_done         <= 0;
                  spc561_phy_pc_w          <= 0;
                end else begin
                  active_thread[(561*4)]   <= 1'b1;
                  active_thread[(561*4)+1] <= 1'b1;
                  active_thread[(561*4)+2] <= 1'b1;
                  active_thread[(561*4)+3] <= 1'b1;
                  spc561_inst_done         <= `ARIANE_CORE561.piton_pc_vld;
                  spc561_phy_pc_w          <= `ARIANE_CORE561.piton_pc;
                end
            end
    

            assign spc562_thread_id = 2'b00;
            assign spc562_rtl_pc = spc562_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(562*4)]   <= 1'b0;
                  active_thread[(562*4)+1] <= 1'b0;
                  active_thread[(562*4)+2] <= 1'b0;
                  active_thread[(562*4)+3] <= 1'b0;
                  spc562_inst_done         <= 0;
                  spc562_phy_pc_w          <= 0;
                end else begin
                  active_thread[(562*4)]   <= 1'b1;
                  active_thread[(562*4)+1] <= 1'b1;
                  active_thread[(562*4)+2] <= 1'b1;
                  active_thread[(562*4)+3] <= 1'b1;
                  spc562_inst_done         <= `ARIANE_CORE562.piton_pc_vld;
                  spc562_phy_pc_w          <= `ARIANE_CORE562.piton_pc;
                end
            end
    

            assign spc563_thread_id = 2'b00;
            assign spc563_rtl_pc = spc563_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(563*4)]   <= 1'b0;
                  active_thread[(563*4)+1] <= 1'b0;
                  active_thread[(563*4)+2] <= 1'b0;
                  active_thread[(563*4)+3] <= 1'b0;
                  spc563_inst_done         <= 0;
                  spc563_phy_pc_w          <= 0;
                end else begin
                  active_thread[(563*4)]   <= 1'b1;
                  active_thread[(563*4)+1] <= 1'b1;
                  active_thread[(563*4)+2] <= 1'b1;
                  active_thread[(563*4)+3] <= 1'b1;
                  spc563_inst_done         <= `ARIANE_CORE563.piton_pc_vld;
                  spc563_phy_pc_w          <= `ARIANE_CORE563.piton_pc;
                end
            end
    

            assign spc564_thread_id = 2'b00;
            assign spc564_rtl_pc = spc564_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(564*4)]   <= 1'b0;
                  active_thread[(564*4)+1] <= 1'b0;
                  active_thread[(564*4)+2] <= 1'b0;
                  active_thread[(564*4)+3] <= 1'b0;
                  spc564_inst_done         <= 0;
                  spc564_phy_pc_w          <= 0;
                end else begin
                  active_thread[(564*4)]   <= 1'b1;
                  active_thread[(564*4)+1] <= 1'b1;
                  active_thread[(564*4)+2] <= 1'b1;
                  active_thread[(564*4)+3] <= 1'b1;
                  spc564_inst_done         <= `ARIANE_CORE564.piton_pc_vld;
                  spc564_phy_pc_w          <= `ARIANE_CORE564.piton_pc;
                end
            end
    

            assign spc565_thread_id = 2'b00;
            assign spc565_rtl_pc = spc565_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(565*4)]   <= 1'b0;
                  active_thread[(565*4)+1] <= 1'b0;
                  active_thread[(565*4)+2] <= 1'b0;
                  active_thread[(565*4)+3] <= 1'b0;
                  spc565_inst_done         <= 0;
                  spc565_phy_pc_w          <= 0;
                end else begin
                  active_thread[(565*4)]   <= 1'b1;
                  active_thread[(565*4)+1] <= 1'b1;
                  active_thread[(565*4)+2] <= 1'b1;
                  active_thread[(565*4)+3] <= 1'b1;
                  spc565_inst_done         <= `ARIANE_CORE565.piton_pc_vld;
                  spc565_phy_pc_w          <= `ARIANE_CORE565.piton_pc;
                end
            end
    

            assign spc566_thread_id = 2'b00;
            assign spc566_rtl_pc = spc566_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(566*4)]   <= 1'b0;
                  active_thread[(566*4)+1] <= 1'b0;
                  active_thread[(566*4)+2] <= 1'b0;
                  active_thread[(566*4)+3] <= 1'b0;
                  spc566_inst_done         <= 0;
                  spc566_phy_pc_w          <= 0;
                end else begin
                  active_thread[(566*4)]   <= 1'b1;
                  active_thread[(566*4)+1] <= 1'b1;
                  active_thread[(566*4)+2] <= 1'b1;
                  active_thread[(566*4)+3] <= 1'b1;
                  spc566_inst_done         <= `ARIANE_CORE566.piton_pc_vld;
                  spc566_phy_pc_w          <= `ARIANE_CORE566.piton_pc;
                end
            end
    

            assign spc567_thread_id = 2'b00;
            assign spc567_rtl_pc = spc567_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(567*4)]   <= 1'b0;
                  active_thread[(567*4)+1] <= 1'b0;
                  active_thread[(567*4)+2] <= 1'b0;
                  active_thread[(567*4)+3] <= 1'b0;
                  spc567_inst_done         <= 0;
                  spc567_phy_pc_w          <= 0;
                end else begin
                  active_thread[(567*4)]   <= 1'b1;
                  active_thread[(567*4)+1] <= 1'b1;
                  active_thread[(567*4)+2] <= 1'b1;
                  active_thread[(567*4)+3] <= 1'b1;
                  spc567_inst_done         <= `ARIANE_CORE567.piton_pc_vld;
                  spc567_phy_pc_w          <= `ARIANE_CORE567.piton_pc;
                end
            end
    

            assign spc568_thread_id = 2'b00;
            assign spc568_rtl_pc = spc568_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(568*4)]   <= 1'b0;
                  active_thread[(568*4)+1] <= 1'b0;
                  active_thread[(568*4)+2] <= 1'b0;
                  active_thread[(568*4)+3] <= 1'b0;
                  spc568_inst_done         <= 0;
                  spc568_phy_pc_w          <= 0;
                end else begin
                  active_thread[(568*4)]   <= 1'b1;
                  active_thread[(568*4)+1] <= 1'b1;
                  active_thread[(568*4)+2] <= 1'b1;
                  active_thread[(568*4)+3] <= 1'b1;
                  spc568_inst_done         <= `ARIANE_CORE568.piton_pc_vld;
                  spc568_phy_pc_w          <= `ARIANE_CORE568.piton_pc;
                end
            end
    

            assign spc569_thread_id = 2'b00;
            assign spc569_rtl_pc = spc569_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(569*4)]   <= 1'b0;
                  active_thread[(569*4)+1] <= 1'b0;
                  active_thread[(569*4)+2] <= 1'b0;
                  active_thread[(569*4)+3] <= 1'b0;
                  spc569_inst_done         <= 0;
                  spc569_phy_pc_w          <= 0;
                end else begin
                  active_thread[(569*4)]   <= 1'b1;
                  active_thread[(569*4)+1] <= 1'b1;
                  active_thread[(569*4)+2] <= 1'b1;
                  active_thread[(569*4)+3] <= 1'b1;
                  spc569_inst_done         <= `ARIANE_CORE569.piton_pc_vld;
                  spc569_phy_pc_w          <= `ARIANE_CORE569.piton_pc;
                end
            end
    

            assign spc570_thread_id = 2'b00;
            assign spc570_rtl_pc = spc570_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(570*4)]   <= 1'b0;
                  active_thread[(570*4)+1] <= 1'b0;
                  active_thread[(570*4)+2] <= 1'b0;
                  active_thread[(570*4)+3] <= 1'b0;
                  spc570_inst_done         <= 0;
                  spc570_phy_pc_w          <= 0;
                end else begin
                  active_thread[(570*4)]   <= 1'b1;
                  active_thread[(570*4)+1] <= 1'b1;
                  active_thread[(570*4)+2] <= 1'b1;
                  active_thread[(570*4)+3] <= 1'b1;
                  spc570_inst_done         <= `ARIANE_CORE570.piton_pc_vld;
                  spc570_phy_pc_w          <= `ARIANE_CORE570.piton_pc;
                end
            end
    

            assign spc571_thread_id = 2'b00;
            assign spc571_rtl_pc = spc571_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(571*4)]   <= 1'b0;
                  active_thread[(571*4)+1] <= 1'b0;
                  active_thread[(571*4)+2] <= 1'b0;
                  active_thread[(571*4)+3] <= 1'b0;
                  spc571_inst_done         <= 0;
                  spc571_phy_pc_w          <= 0;
                end else begin
                  active_thread[(571*4)]   <= 1'b1;
                  active_thread[(571*4)+1] <= 1'b1;
                  active_thread[(571*4)+2] <= 1'b1;
                  active_thread[(571*4)+3] <= 1'b1;
                  spc571_inst_done         <= `ARIANE_CORE571.piton_pc_vld;
                  spc571_phy_pc_w          <= `ARIANE_CORE571.piton_pc;
                end
            end
    

            assign spc572_thread_id = 2'b00;
            assign spc572_rtl_pc = spc572_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(572*4)]   <= 1'b0;
                  active_thread[(572*4)+1] <= 1'b0;
                  active_thread[(572*4)+2] <= 1'b0;
                  active_thread[(572*4)+3] <= 1'b0;
                  spc572_inst_done         <= 0;
                  spc572_phy_pc_w          <= 0;
                end else begin
                  active_thread[(572*4)]   <= 1'b1;
                  active_thread[(572*4)+1] <= 1'b1;
                  active_thread[(572*4)+2] <= 1'b1;
                  active_thread[(572*4)+3] <= 1'b1;
                  spc572_inst_done         <= `ARIANE_CORE572.piton_pc_vld;
                  spc572_phy_pc_w          <= `ARIANE_CORE572.piton_pc;
                end
            end
    

            assign spc573_thread_id = 2'b00;
            assign spc573_rtl_pc = spc573_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(573*4)]   <= 1'b0;
                  active_thread[(573*4)+1] <= 1'b0;
                  active_thread[(573*4)+2] <= 1'b0;
                  active_thread[(573*4)+3] <= 1'b0;
                  spc573_inst_done         <= 0;
                  spc573_phy_pc_w          <= 0;
                end else begin
                  active_thread[(573*4)]   <= 1'b1;
                  active_thread[(573*4)+1] <= 1'b1;
                  active_thread[(573*4)+2] <= 1'b1;
                  active_thread[(573*4)+3] <= 1'b1;
                  spc573_inst_done         <= `ARIANE_CORE573.piton_pc_vld;
                  spc573_phy_pc_w          <= `ARIANE_CORE573.piton_pc;
                end
            end
    

            assign spc574_thread_id = 2'b00;
            assign spc574_rtl_pc = spc574_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(574*4)]   <= 1'b0;
                  active_thread[(574*4)+1] <= 1'b0;
                  active_thread[(574*4)+2] <= 1'b0;
                  active_thread[(574*4)+3] <= 1'b0;
                  spc574_inst_done         <= 0;
                  spc574_phy_pc_w          <= 0;
                end else begin
                  active_thread[(574*4)]   <= 1'b1;
                  active_thread[(574*4)+1] <= 1'b1;
                  active_thread[(574*4)+2] <= 1'b1;
                  active_thread[(574*4)+3] <= 1'b1;
                  spc574_inst_done         <= `ARIANE_CORE574.piton_pc_vld;
                  spc574_phy_pc_w          <= `ARIANE_CORE574.piton_pc;
                end
            end
    

            assign spc575_thread_id = 2'b00;
            assign spc575_rtl_pc = spc575_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(575*4)]   <= 1'b0;
                  active_thread[(575*4)+1] <= 1'b0;
                  active_thread[(575*4)+2] <= 1'b0;
                  active_thread[(575*4)+3] <= 1'b0;
                  spc575_inst_done         <= 0;
                  spc575_phy_pc_w          <= 0;
                end else begin
                  active_thread[(575*4)]   <= 1'b1;
                  active_thread[(575*4)+1] <= 1'b1;
                  active_thread[(575*4)+2] <= 1'b1;
                  active_thread[(575*4)+3] <= 1'b1;
                  spc575_inst_done         <= `ARIANE_CORE575.piton_pc_vld;
                  spc575_phy_pc_w          <= `ARIANE_CORE575.piton_pc;
                end
            end
    

            assign spc576_thread_id = 2'b00;
            assign spc576_rtl_pc = spc576_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(576*4)]   <= 1'b0;
                  active_thread[(576*4)+1] <= 1'b0;
                  active_thread[(576*4)+2] <= 1'b0;
                  active_thread[(576*4)+3] <= 1'b0;
                  spc576_inst_done         <= 0;
                  spc576_phy_pc_w          <= 0;
                end else begin
                  active_thread[(576*4)]   <= 1'b1;
                  active_thread[(576*4)+1] <= 1'b1;
                  active_thread[(576*4)+2] <= 1'b1;
                  active_thread[(576*4)+3] <= 1'b1;
                  spc576_inst_done         <= `ARIANE_CORE576.piton_pc_vld;
                  spc576_phy_pc_w          <= `ARIANE_CORE576.piton_pc;
                end
            end
    

            assign spc577_thread_id = 2'b00;
            assign spc577_rtl_pc = spc577_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(577*4)]   <= 1'b0;
                  active_thread[(577*4)+1] <= 1'b0;
                  active_thread[(577*4)+2] <= 1'b0;
                  active_thread[(577*4)+3] <= 1'b0;
                  spc577_inst_done         <= 0;
                  spc577_phy_pc_w          <= 0;
                end else begin
                  active_thread[(577*4)]   <= 1'b1;
                  active_thread[(577*4)+1] <= 1'b1;
                  active_thread[(577*4)+2] <= 1'b1;
                  active_thread[(577*4)+3] <= 1'b1;
                  spc577_inst_done         <= `ARIANE_CORE577.piton_pc_vld;
                  spc577_phy_pc_w          <= `ARIANE_CORE577.piton_pc;
                end
            end
    

            assign spc578_thread_id = 2'b00;
            assign spc578_rtl_pc = spc578_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(578*4)]   <= 1'b0;
                  active_thread[(578*4)+1] <= 1'b0;
                  active_thread[(578*4)+2] <= 1'b0;
                  active_thread[(578*4)+3] <= 1'b0;
                  spc578_inst_done         <= 0;
                  spc578_phy_pc_w          <= 0;
                end else begin
                  active_thread[(578*4)]   <= 1'b1;
                  active_thread[(578*4)+1] <= 1'b1;
                  active_thread[(578*4)+2] <= 1'b1;
                  active_thread[(578*4)+3] <= 1'b1;
                  spc578_inst_done         <= `ARIANE_CORE578.piton_pc_vld;
                  spc578_phy_pc_w          <= `ARIANE_CORE578.piton_pc;
                end
            end
    

            assign spc579_thread_id = 2'b00;
            assign spc579_rtl_pc = spc579_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(579*4)]   <= 1'b0;
                  active_thread[(579*4)+1] <= 1'b0;
                  active_thread[(579*4)+2] <= 1'b0;
                  active_thread[(579*4)+3] <= 1'b0;
                  spc579_inst_done         <= 0;
                  spc579_phy_pc_w          <= 0;
                end else begin
                  active_thread[(579*4)]   <= 1'b1;
                  active_thread[(579*4)+1] <= 1'b1;
                  active_thread[(579*4)+2] <= 1'b1;
                  active_thread[(579*4)+3] <= 1'b1;
                  spc579_inst_done         <= `ARIANE_CORE579.piton_pc_vld;
                  spc579_phy_pc_w          <= `ARIANE_CORE579.piton_pc;
                end
            end
    

            assign spc580_thread_id = 2'b00;
            assign spc580_rtl_pc = spc580_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(580*4)]   <= 1'b0;
                  active_thread[(580*4)+1] <= 1'b0;
                  active_thread[(580*4)+2] <= 1'b0;
                  active_thread[(580*4)+3] <= 1'b0;
                  spc580_inst_done         <= 0;
                  spc580_phy_pc_w          <= 0;
                end else begin
                  active_thread[(580*4)]   <= 1'b1;
                  active_thread[(580*4)+1] <= 1'b1;
                  active_thread[(580*4)+2] <= 1'b1;
                  active_thread[(580*4)+3] <= 1'b1;
                  spc580_inst_done         <= `ARIANE_CORE580.piton_pc_vld;
                  spc580_phy_pc_w          <= `ARIANE_CORE580.piton_pc;
                end
            end
    

            assign spc581_thread_id = 2'b00;
            assign spc581_rtl_pc = spc581_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(581*4)]   <= 1'b0;
                  active_thread[(581*4)+1] <= 1'b0;
                  active_thread[(581*4)+2] <= 1'b0;
                  active_thread[(581*4)+3] <= 1'b0;
                  spc581_inst_done         <= 0;
                  spc581_phy_pc_w          <= 0;
                end else begin
                  active_thread[(581*4)]   <= 1'b1;
                  active_thread[(581*4)+1] <= 1'b1;
                  active_thread[(581*4)+2] <= 1'b1;
                  active_thread[(581*4)+3] <= 1'b1;
                  spc581_inst_done         <= `ARIANE_CORE581.piton_pc_vld;
                  spc581_phy_pc_w          <= `ARIANE_CORE581.piton_pc;
                end
            end
    

            assign spc582_thread_id = 2'b00;
            assign spc582_rtl_pc = spc582_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(582*4)]   <= 1'b0;
                  active_thread[(582*4)+1] <= 1'b0;
                  active_thread[(582*4)+2] <= 1'b0;
                  active_thread[(582*4)+3] <= 1'b0;
                  spc582_inst_done         <= 0;
                  spc582_phy_pc_w          <= 0;
                end else begin
                  active_thread[(582*4)]   <= 1'b1;
                  active_thread[(582*4)+1] <= 1'b1;
                  active_thread[(582*4)+2] <= 1'b1;
                  active_thread[(582*4)+3] <= 1'b1;
                  spc582_inst_done         <= `ARIANE_CORE582.piton_pc_vld;
                  spc582_phy_pc_w          <= `ARIANE_CORE582.piton_pc;
                end
            end
    

            assign spc583_thread_id = 2'b00;
            assign spc583_rtl_pc = spc583_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(583*4)]   <= 1'b0;
                  active_thread[(583*4)+1] <= 1'b0;
                  active_thread[(583*4)+2] <= 1'b0;
                  active_thread[(583*4)+3] <= 1'b0;
                  spc583_inst_done         <= 0;
                  spc583_phy_pc_w          <= 0;
                end else begin
                  active_thread[(583*4)]   <= 1'b1;
                  active_thread[(583*4)+1] <= 1'b1;
                  active_thread[(583*4)+2] <= 1'b1;
                  active_thread[(583*4)+3] <= 1'b1;
                  spc583_inst_done         <= `ARIANE_CORE583.piton_pc_vld;
                  spc583_phy_pc_w          <= `ARIANE_CORE583.piton_pc;
                end
            end
    

            assign spc584_thread_id = 2'b00;
            assign spc584_rtl_pc = spc584_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(584*4)]   <= 1'b0;
                  active_thread[(584*4)+1] <= 1'b0;
                  active_thread[(584*4)+2] <= 1'b0;
                  active_thread[(584*4)+3] <= 1'b0;
                  spc584_inst_done         <= 0;
                  spc584_phy_pc_w          <= 0;
                end else begin
                  active_thread[(584*4)]   <= 1'b1;
                  active_thread[(584*4)+1] <= 1'b1;
                  active_thread[(584*4)+2] <= 1'b1;
                  active_thread[(584*4)+3] <= 1'b1;
                  spc584_inst_done         <= `ARIANE_CORE584.piton_pc_vld;
                  spc584_phy_pc_w          <= `ARIANE_CORE584.piton_pc;
                end
            end
    

            assign spc585_thread_id = 2'b00;
            assign spc585_rtl_pc = spc585_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(585*4)]   <= 1'b0;
                  active_thread[(585*4)+1] <= 1'b0;
                  active_thread[(585*4)+2] <= 1'b0;
                  active_thread[(585*4)+3] <= 1'b0;
                  spc585_inst_done         <= 0;
                  spc585_phy_pc_w          <= 0;
                end else begin
                  active_thread[(585*4)]   <= 1'b1;
                  active_thread[(585*4)+1] <= 1'b1;
                  active_thread[(585*4)+2] <= 1'b1;
                  active_thread[(585*4)+3] <= 1'b1;
                  spc585_inst_done         <= `ARIANE_CORE585.piton_pc_vld;
                  spc585_phy_pc_w          <= `ARIANE_CORE585.piton_pc;
                end
            end
    

            assign spc586_thread_id = 2'b00;
            assign spc586_rtl_pc = spc586_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(586*4)]   <= 1'b0;
                  active_thread[(586*4)+1] <= 1'b0;
                  active_thread[(586*4)+2] <= 1'b0;
                  active_thread[(586*4)+3] <= 1'b0;
                  spc586_inst_done         <= 0;
                  spc586_phy_pc_w          <= 0;
                end else begin
                  active_thread[(586*4)]   <= 1'b1;
                  active_thread[(586*4)+1] <= 1'b1;
                  active_thread[(586*4)+2] <= 1'b1;
                  active_thread[(586*4)+3] <= 1'b1;
                  spc586_inst_done         <= `ARIANE_CORE586.piton_pc_vld;
                  spc586_phy_pc_w          <= `ARIANE_CORE586.piton_pc;
                end
            end
    

            assign spc587_thread_id = 2'b00;
            assign spc587_rtl_pc = spc587_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(587*4)]   <= 1'b0;
                  active_thread[(587*4)+1] <= 1'b0;
                  active_thread[(587*4)+2] <= 1'b0;
                  active_thread[(587*4)+3] <= 1'b0;
                  spc587_inst_done         <= 0;
                  spc587_phy_pc_w          <= 0;
                end else begin
                  active_thread[(587*4)]   <= 1'b1;
                  active_thread[(587*4)+1] <= 1'b1;
                  active_thread[(587*4)+2] <= 1'b1;
                  active_thread[(587*4)+3] <= 1'b1;
                  spc587_inst_done         <= `ARIANE_CORE587.piton_pc_vld;
                  spc587_phy_pc_w          <= `ARIANE_CORE587.piton_pc;
                end
            end
    

            assign spc588_thread_id = 2'b00;
            assign spc588_rtl_pc = spc588_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(588*4)]   <= 1'b0;
                  active_thread[(588*4)+1] <= 1'b0;
                  active_thread[(588*4)+2] <= 1'b0;
                  active_thread[(588*4)+3] <= 1'b0;
                  spc588_inst_done         <= 0;
                  spc588_phy_pc_w          <= 0;
                end else begin
                  active_thread[(588*4)]   <= 1'b1;
                  active_thread[(588*4)+1] <= 1'b1;
                  active_thread[(588*4)+2] <= 1'b1;
                  active_thread[(588*4)+3] <= 1'b1;
                  spc588_inst_done         <= `ARIANE_CORE588.piton_pc_vld;
                  spc588_phy_pc_w          <= `ARIANE_CORE588.piton_pc;
                end
            end
    

            assign spc589_thread_id = 2'b00;
            assign spc589_rtl_pc = spc589_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(589*4)]   <= 1'b0;
                  active_thread[(589*4)+1] <= 1'b0;
                  active_thread[(589*4)+2] <= 1'b0;
                  active_thread[(589*4)+3] <= 1'b0;
                  spc589_inst_done         <= 0;
                  spc589_phy_pc_w          <= 0;
                end else begin
                  active_thread[(589*4)]   <= 1'b1;
                  active_thread[(589*4)+1] <= 1'b1;
                  active_thread[(589*4)+2] <= 1'b1;
                  active_thread[(589*4)+3] <= 1'b1;
                  spc589_inst_done         <= `ARIANE_CORE589.piton_pc_vld;
                  spc589_phy_pc_w          <= `ARIANE_CORE589.piton_pc;
                end
            end
    

            assign spc590_thread_id = 2'b00;
            assign spc590_rtl_pc = spc590_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(590*4)]   <= 1'b0;
                  active_thread[(590*4)+1] <= 1'b0;
                  active_thread[(590*4)+2] <= 1'b0;
                  active_thread[(590*4)+3] <= 1'b0;
                  spc590_inst_done         <= 0;
                  spc590_phy_pc_w          <= 0;
                end else begin
                  active_thread[(590*4)]   <= 1'b1;
                  active_thread[(590*4)+1] <= 1'b1;
                  active_thread[(590*4)+2] <= 1'b1;
                  active_thread[(590*4)+3] <= 1'b1;
                  spc590_inst_done         <= `ARIANE_CORE590.piton_pc_vld;
                  spc590_phy_pc_w          <= `ARIANE_CORE590.piton_pc;
                end
            end
    

            assign spc591_thread_id = 2'b00;
            assign spc591_rtl_pc = spc591_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(591*4)]   <= 1'b0;
                  active_thread[(591*4)+1] <= 1'b0;
                  active_thread[(591*4)+2] <= 1'b0;
                  active_thread[(591*4)+3] <= 1'b0;
                  spc591_inst_done         <= 0;
                  spc591_phy_pc_w          <= 0;
                end else begin
                  active_thread[(591*4)]   <= 1'b1;
                  active_thread[(591*4)+1] <= 1'b1;
                  active_thread[(591*4)+2] <= 1'b1;
                  active_thread[(591*4)+3] <= 1'b1;
                  spc591_inst_done         <= `ARIANE_CORE591.piton_pc_vld;
                  spc591_phy_pc_w          <= `ARIANE_CORE591.piton_pc;
                end
            end
    

            assign spc592_thread_id = 2'b00;
            assign spc592_rtl_pc = spc592_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(592*4)]   <= 1'b0;
                  active_thread[(592*4)+1] <= 1'b0;
                  active_thread[(592*4)+2] <= 1'b0;
                  active_thread[(592*4)+3] <= 1'b0;
                  spc592_inst_done         <= 0;
                  spc592_phy_pc_w          <= 0;
                end else begin
                  active_thread[(592*4)]   <= 1'b1;
                  active_thread[(592*4)+1] <= 1'b1;
                  active_thread[(592*4)+2] <= 1'b1;
                  active_thread[(592*4)+3] <= 1'b1;
                  spc592_inst_done         <= `ARIANE_CORE592.piton_pc_vld;
                  spc592_phy_pc_w          <= `ARIANE_CORE592.piton_pc;
                end
            end
    

            assign spc593_thread_id = 2'b00;
            assign spc593_rtl_pc = spc593_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(593*4)]   <= 1'b0;
                  active_thread[(593*4)+1] <= 1'b0;
                  active_thread[(593*4)+2] <= 1'b0;
                  active_thread[(593*4)+3] <= 1'b0;
                  spc593_inst_done         <= 0;
                  spc593_phy_pc_w          <= 0;
                end else begin
                  active_thread[(593*4)]   <= 1'b1;
                  active_thread[(593*4)+1] <= 1'b1;
                  active_thread[(593*4)+2] <= 1'b1;
                  active_thread[(593*4)+3] <= 1'b1;
                  spc593_inst_done         <= `ARIANE_CORE593.piton_pc_vld;
                  spc593_phy_pc_w          <= `ARIANE_CORE593.piton_pc;
                end
            end
    

            assign spc594_thread_id = 2'b00;
            assign spc594_rtl_pc = spc594_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(594*4)]   <= 1'b0;
                  active_thread[(594*4)+1] <= 1'b0;
                  active_thread[(594*4)+2] <= 1'b0;
                  active_thread[(594*4)+3] <= 1'b0;
                  spc594_inst_done         <= 0;
                  spc594_phy_pc_w          <= 0;
                end else begin
                  active_thread[(594*4)]   <= 1'b1;
                  active_thread[(594*4)+1] <= 1'b1;
                  active_thread[(594*4)+2] <= 1'b1;
                  active_thread[(594*4)+3] <= 1'b1;
                  spc594_inst_done         <= `ARIANE_CORE594.piton_pc_vld;
                  spc594_phy_pc_w          <= `ARIANE_CORE594.piton_pc;
                end
            end
    

            assign spc595_thread_id = 2'b00;
            assign spc595_rtl_pc = spc595_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(595*4)]   <= 1'b0;
                  active_thread[(595*4)+1] <= 1'b0;
                  active_thread[(595*4)+2] <= 1'b0;
                  active_thread[(595*4)+3] <= 1'b0;
                  spc595_inst_done         <= 0;
                  spc595_phy_pc_w          <= 0;
                end else begin
                  active_thread[(595*4)]   <= 1'b1;
                  active_thread[(595*4)+1] <= 1'b1;
                  active_thread[(595*4)+2] <= 1'b1;
                  active_thread[(595*4)+3] <= 1'b1;
                  spc595_inst_done         <= `ARIANE_CORE595.piton_pc_vld;
                  spc595_phy_pc_w          <= `ARIANE_CORE595.piton_pc;
                end
            end
    

            assign spc596_thread_id = 2'b00;
            assign spc596_rtl_pc = spc596_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(596*4)]   <= 1'b0;
                  active_thread[(596*4)+1] <= 1'b0;
                  active_thread[(596*4)+2] <= 1'b0;
                  active_thread[(596*4)+3] <= 1'b0;
                  spc596_inst_done         <= 0;
                  spc596_phy_pc_w          <= 0;
                end else begin
                  active_thread[(596*4)]   <= 1'b1;
                  active_thread[(596*4)+1] <= 1'b1;
                  active_thread[(596*4)+2] <= 1'b1;
                  active_thread[(596*4)+3] <= 1'b1;
                  spc596_inst_done         <= `ARIANE_CORE596.piton_pc_vld;
                  spc596_phy_pc_w          <= `ARIANE_CORE596.piton_pc;
                end
            end
    

            assign spc597_thread_id = 2'b00;
            assign spc597_rtl_pc = spc597_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(597*4)]   <= 1'b0;
                  active_thread[(597*4)+1] <= 1'b0;
                  active_thread[(597*4)+2] <= 1'b0;
                  active_thread[(597*4)+3] <= 1'b0;
                  spc597_inst_done         <= 0;
                  spc597_phy_pc_w          <= 0;
                end else begin
                  active_thread[(597*4)]   <= 1'b1;
                  active_thread[(597*4)+1] <= 1'b1;
                  active_thread[(597*4)+2] <= 1'b1;
                  active_thread[(597*4)+3] <= 1'b1;
                  spc597_inst_done         <= `ARIANE_CORE597.piton_pc_vld;
                  spc597_phy_pc_w          <= `ARIANE_CORE597.piton_pc;
                end
            end
    

            assign spc598_thread_id = 2'b00;
            assign spc598_rtl_pc = spc598_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(598*4)]   <= 1'b0;
                  active_thread[(598*4)+1] <= 1'b0;
                  active_thread[(598*4)+2] <= 1'b0;
                  active_thread[(598*4)+3] <= 1'b0;
                  spc598_inst_done         <= 0;
                  spc598_phy_pc_w          <= 0;
                end else begin
                  active_thread[(598*4)]   <= 1'b1;
                  active_thread[(598*4)+1] <= 1'b1;
                  active_thread[(598*4)+2] <= 1'b1;
                  active_thread[(598*4)+3] <= 1'b1;
                  spc598_inst_done         <= `ARIANE_CORE598.piton_pc_vld;
                  spc598_phy_pc_w          <= `ARIANE_CORE598.piton_pc;
                end
            end
    

            assign spc599_thread_id = 2'b00;
            assign spc599_rtl_pc = spc599_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(599*4)]   <= 1'b0;
                  active_thread[(599*4)+1] <= 1'b0;
                  active_thread[(599*4)+2] <= 1'b0;
                  active_thread[(599*4)+3] <= 1'b0;
                  spc599_inst_done         <= 0;
                  spc599_phy_pc_w          <= 0;
                end else begin
                  active_thread[(599*4)]   <= 1'b1;
                  active_thread[(599*4)+1] <= 1'b1;
                  active_thread[(599*4)+2] <= 1'b1;
                  active_thread[(599*4)+3] <= 1'b1;
                  spc599_inst_done         <= `ARIANE_CORE599.piton_pc_vld;
                  spc599_phy_pc_w          <= `ARIANE_CORE599.piton_pc;
                end
            end
    

            assign spc600_thread_id = 2'b00;
            assign spc600_rtl_pc = spc600_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(600*4)]   <= 1'b0;
                  active_thread[(600*4)+1] <= 1'b0;
                  active_thread[(600*4)+2] <= 1'b0;
                  active_thread[(600*4)+3] <= 1'b0;
                  spc600_inst_done         <= 0;
                  spc600_phy_pc_w          <= 0;
                end else begin
                  active_thread[(600*4)]   <= 1'b1;
                  active_thread[(600*4)+1] <= 1'b1;
                  active_thread[(600*4)+2] <= 1'b1;
                  active_thread[(600*4)+3] <= 1'b1;
                  spc600_inst_done         <= `ARIANE_CORE600.piton_pc_vld;
                  spc600_phy_pc_w          <= `ARIANE_CORE600.piton_pc;
                end
            end
    

            assign spc601_thread_id = 2'b00;
            assign spc601_rtl_pc = spc601_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(601*4)]   <= 1'b0;
                  active_thread[(601*4)+1] <= 1'b0;
                  active_thread[(601*4)+2] <= 1'b0;
                  active_thread[(601*4)+3] <= 1'b0;
                  spc601_inst_done         <= 0;
                  spc601_phy_pc_w          <= 0;
                end else begin
                  active_thread[(601*4)]   <= 1'b1;
                  active_thread[(601*4)+1] <= 1'b1;
                  active_thread[(601*4)+2] <= 1'b1;
                  active_thread[(601*4)+3] <= 1'b1;
                  spc601_inst_done         <= `ARIANE_CORE601.piton_pc_vld;
                  spc601_phy_pc_w          <= `ARIANE_CORE601.piton_pc;
                end
            end
    

            assign spc602_thread_id = 2'b00;
            assign spc602_rtl_pc = spc602_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(602*4)]   <= 1'b0;
                  active_thread[(602*4)+1] <= 1'b0;
                  active_thread[(602*4)+2] <= 1'b0;
                  active_thread[(602*4)+3] <= 1'b0;
                  spc602_inst_done         <= 0;
                  spc602_phy_pc_w          <= 0;
                end else begin
                  active_thread[(602*4)]   <= 1'b1;
                  active_thread[(602*4)+1] <= 1'b1;
                  active_thread[(602*4)+2] <= 1'b1;
                  active_thread[(602*4)+3] <= 1'b1;
                  spc602_inst_done         <= `ARIANE_CORE602.piton_pc_vld;
                  spc602_phy_pc_w          <= `ARIANE_CORE602.piton_pc;
                end
            end
    

            assign spc603_thread_id = 2'b00;
            assign spc603_rtl_pc = spc603_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(603*4)]   <= 1'b0;
                  active_thread[(603*4)+1] <= 1'b0;
                  active_thread[(603*4)+2] <= 1'b0;
                  active_thread[(603*4)+3] <= 1'b0;
                  spc603_inst_done         <= 0;
                  spc603_phy_pc_w          <= 0;
                end else begin
                  active_thread[(603*4)]   <= 1'b1;
                  active_thread[(603*4)+1] <= 1'b1;
                  active_thread[(603*4)+2] <= 1'b1;
                  active_thread[(603*4)+3] <= 1'b1;
                  spc603_inst_done         <= `ARIANE_CORE603.piton_pc_vld;
                  spc603_phy_pc_w          <= `ARIANE_CORE603.piton_pc;
                end
            end
    

            assign spc604_thread_id = 2'b00;
            assign spc604_rtl_pc = spc604_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(604*4)]   <= 1'b0;
                  active_thread[(604*4)+1] <= 1'b0;
                  active_thread[(604*4)+2] <= 1'b0;
                  active_thread[(604*4)+3] <= 1'b0;
                  spc604_inst_done         <= 0;
                  spc604_phy_pc_w          <= 0;
                end else begin
                  active_thread[(604*4)]   <= 1'b1;
                  active_thread[(604*4)+1] <= 1'b1;
                  active_thread[(604*4)+2] <= 1'b1;
                  active_thread[(604*4)+3] <= 1'b1;
                  spc604_inst_done         <= `ARIANE_CORE604.piton_pc_vld;
                  spc604_phy_pc_w          <= `ARIANE_CORE604.piton_pc;
                end
            end
    

            assign spc605_thread_id = 2'b00;
            assign spc605_rtl_pc = spc605_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(605*4)]   <= 1'b0;
                  active_thread[(605*4)+1] <= 1'b0;
                  active_thread[(605*4)+2] <= 1'b0;
                  active_thread[(605*4)+3] <= 1'b0;
                  spc605_inst_done         <= 0;
                  spc605_phy_pc_w          <= 0;
                end else begin
                  active_thread[(605*4)]   <= 1'b1;
                  active_thread[(605*4)+1] <= 1'b1;
                  active_thread[(605*4)+2] <= 1'b1;
                  active_thread[(605*4)+3] <= 1'b1;
                  spc605_inst_done         <= `ARIANE_CORE605.piton_pc_vld;
                  spc605_phy_pc_w          <= `ARIANE_CORE605.piton_pc;
                end
            end
    

            assign spc606_thread_id = 2'b00;
            assign spc606_rtl_pc = spc606_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(606*4)]   <= 1'b0;
                  active_thread[(606*4)+1] <= 1'b0;
                  active_thread[(606*4)+2] <= 1'b0;
                  active_thread[(606*4)+3] <= 1'b0;
                  spc606_inst_done         <= 0;
                  spc606_phy_pc_w          <= 0;
                end else begin
                  active_thread[(606*4)]   <= 1'b1;
                  active_thread[(606*4)+1] <= 1'b1;
                  active_thread[(606*4)+2] <= 1'b1;
                  active_thread[(606*4)+3] <= 1'b1;
                  spc606_inst_done         <= `ARIANE_CORE606.piton_pc_vld;
                  spc606_phy_pc_w          <= `ARIANE_CORE606.piton_pc;
                end
            end
    

            assign spc607_thread_id = 2'b00;
            assign spc607_rtl_pc = spc607_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(607*4)]   <= 1'b0;
                  active_thread[(607*4)+1] <= 1'b0;
                  active_thread[(607*4)+2] <= 1'b0;
                  active_thread[(607*4)+3] <= 1'b0;
                  spc607_inst_done         <= 0;
                  spc607_phy_pc_w          <= 0;
                end else begin
                  active_thread[(607*4)]   <= 1'b1;
                  active_thread[(607*4)+1] <= 1'b1;
                  active_thread[(607*4)+2] <= 1'b1;
                  active_thread[(607*4)+3] <= 1'b1;
                  spc607_inst_done         <= `ARIANE_CORE607.piton_pc_vld;
                  spc607_phy_pc_w          <= `ARIANE_CORE607.piton_pc;
                end
            end
    

            assign spc608_thread_id = 2'b00;
            assign spc608_rtl_pc = spc608_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(608*4)]   <= 1'b0;
                  active_thread[(608*4)+1] <= 1'b0;
                  active_thread[(608*4)+2] <= 1'b0;
                  active_thread[(608*4)+3] <= 1'b0;
                  spc608_inst_done         <= 0;
                  spc608_phy_pc_w          <= 0;
                end else begin
                  active_thread[(608*4)]   <= 1'b1;
                  active_thread[(608*4)+1] <= 1'b1;
                  active_thread[(608*4)+2] <= 1'b1;
                  active_thread[(608*4)+3] <= 1'b1;
                  spc608_inst_done         <= `ARIANE_CORE608.piton_pc_vld;
                  spc608_phy_pc_w          <= `ARIANE_CORE608.piton_pc;
                end
            end
    

            assign spc609_thread_id = 2'b00;
            assign spc609_rtl_pc = spc609_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(609*4)]   <= 1'b0;
                  active_thread[(609*4)+1] <= 1'b0;
                  active_thread[(609*4)+2] <= 1'b0;
                  active_thread[(609*4)+3] <= 1'b0;
                  spc609_inst_done         <= 0;
                  spc609_phy_pc_w          <= 0;
                end else begin
                  active_thread[(609*4)]   <= 1'b1;
                  active_thread[(609*4)+1] <= 1'b1;
                  active_thread[(609*4)+2] <= 1'b1;
                  active_thread[(609*4)+3] <= 1'b1;
                  spc609_inst_done         <= `ARIANE_CORE609.piton_pc_vld;
                  spc609_phy_pc_w          <= `ARIANE_CORE609.piton_pc;
                end
            end
    

            assign spc610_thread_id = 2'b00;
            assign spc610_rtl_pc = spc610_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(610*4)]   <= 1'b0;
                  active_thread[(610*4)+1] <= 1'b0;
                  active_thread[(610*4)+2] <= 1'b0;
                  active_thread[(610*4)+3] <= 1'b0;
                  spc610_inst_done         <= 0;
                  spc610_phy_pc_w          <= 0;
                end else begin
                  active_thread[(610*4)]   <= 1'b1;
                  active_thread[(610*4)+1] <= 1'b1;
                  active_thread[(610*4)+2] <= 1'b1;
                  active_thread[(610*4)+3] <= 1'b1;
                  spc610_inst_done         <= `ARIANE_CORE610.piton_pc_vld;
                  spc610_phy_pc_w          <= `ARIANE_CORE610.piton_pc;
                end
            end
    

            assign spc611_thread_id = 2'b00;
            assign spc611_rtl_pc = spc611_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(611*4)]   <= 1'b0;
                  active_thread[(611*4)+1] <= 1'b0;
                  active_thread[(611*4)+2] <= 1'b0;
                  active_thread[(611*4)+3] <= 1'b0;
                  spc611_inst_done         <= 0;
                  spc611_phy_pc_w          <= 0;
                end else begin
                  active_thread[(611*4)]   <= 1'b1;
                  active_thread[(611*4)+1] <= 1'b1;
                  active_thread[(611*4)+2] <= 1'b1;
                  active_thread[(611*4)+3] <= 1'b1;
                  spc611_inst_done         <= `ARIANE_CORE611.piton_pc_vld;
                  spc611_phy_pc_w          <= `ARIANE_CORE611.piton_pc;
                end
            end
    

            assign spc612_thread_id = 2'b00;
            assign spc612_rtl_pc = spc612_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(612*4)]   <= 1'b0;
                  active_thread[(612*4)+1] <= 1'b0;
                  active_thread[(612*4)+2] <= 1'b0;
                  active_thread[(612*4)+3] <= 1'b0;
                  spc612_inst_done         <= 0;
                  spc612_phy_pc_w          <= 0;
                end else begin
                  active_thread[(612*4)]   <= 1'b1;
                  active_thread[(612*4)+1] <= 1'b1;
                  active_thread[(612*4)+2] <= 1'b1;
                  active_thread[(612*4)+3] <= 1'b1;
                  spc612_inst_done         <= `ARIANE_CORE612.piton_pc_vld;
                  spc612_phy_pc_w          <= `ARIANE_CORE612.piton_pc;
                end
            end
    

            assign spc613_thread_id = 2'b00;
            assign spc613_rtl_pc = spc613_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(613*4)]   <= 1'b0;
                  active_thread[(613*4)+1] <= 1'b0;
                  active_thread[(613*4)+2] <= 1'b0;
                  active_thread[(613*4)+3] <= 1'b0;
                  spc613_inst_done         <= 0;
                  spc613_phy_pc_w          <= 0;
                end else begin
                  active_thread[(613*4)]   <= 1'b1;
                  active_thread[(613*4)+1] <= 1'b1;
                  active_thread[(613*4)+2] <= 1'b1;
                  active_thread[(613*4)+3] <= 1'b1;
                  spc613_inst_done         <= `ARIANE_CORE613.piton_pc_vld;
                  spc613_phy_pc_w          <= `ARIANE_CORE613.piton_pc;
                end
            end
    

            assign spc614_thread_id = 2'b00;
            assign spc614_rtl_pc = spc614_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(614*4)]   <= 1'b0;
                  active_thread[(614*4)+1] <= 1'b0;
                  active_thread[(614*4)+2] <= 1'b0;
                  active_thread[(614*4)+3] <= 1'b0;
                  spc614_inst_done         <= 0;
                  spc614_phy_pc_w          <= 0;
                end else begin
                  active_thread[(614*4)]   <= 1'b1;
                  active_thread[(614*4)+1] <= 1'b1;
                  active_thread[(614*4)+2] <= 1'b1;
                  active_thread[(614*4)+3] <= 1'b1;
                  spc614_inst_done         <= `ARIANE_CORE614.piton_pc_vld;
                  spc614_phy_pc_w          <= `ARIANE_CORE614.piton_pc;
                end
            end
    

            assign spc615_thread_id = 2'b00;
            assign spc615_rtl_pc = spc615_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(615*4)]   <= 1'b0;
                  active_thread[(615*4)+1] <= 1'b0;
                  active_thread[(615*4)+2] <= 1'b0;
                  active_thread[(615*4)+3] <= 1'b0;
                  spc615_inst_done         <= 0;
                  spc615_phy_pc_w          <= 0;
                end else begin
                  active_thread[(615*4)]   <= 1'b1;
                  active_thread[(615*4)+1] <= 1'b1;
                  active_thread[(615*4)+2] <= 1'b1;
                  active_thread[(615*4)+3] <= 1'b1;
                  spc615_inst_done         <= `ARIANE_CORE615.piton_pc_vld;
                  spc615_phy_pc_w          <= `ARIANE_CORE615.piton_pc;
                end
            end
    

            assign spc616_thread_id = 2'b00;
            assign spc616_rtl_pc = spc616_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(616*4)]   <= 1'b0;
                  active_thread[(616*4)+1] <= 1'b0;
                  active_thread[(616*4)+2] <= 1'b0;
                  active_thread[(616*4)+3] <= 1'b0;
                  spc616_inst_done         <= 0;
                  spc616_phy_pc_w          <= 0;
                end else begin
                  active_thread[(616*4)]   <= 1'b1;
                  active_thread[(616*4)+1] <= 1'b1;
                  active_thread[(616*4)+2] <= 1'b1;
                  active_thread[(616*4)+3] <= 1'b1;
                  spc616_inst_done         <= `ARIANE_CORE616.piton_pc_vld;
                  spc616_phy_pc_w          <= `ARIANE_CORE616.piton_pc;
                end
            end
    

            assign spc617_thread_id = 2'b00;
            assign spc617_rtl_pc = spc617_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(617*4)]   <= 1'b0;
                  active_thread[(617*4)+1] <= 1'b0;
                  active_thread[(617*4)+2] <= 1'b0;
                  active_thread[(617*4)+3] <= 1'b0;
                  spc617_inst_done         <= 0;
                  spc617_phy_pc_w          <= 0;
                end else begin
                  active_thread[(617*4)]   <= 1'b1;
                  active_thread[(617*4)+1] <= 1'b1;
                  active_thread[(617*4)+2] <= 1'b1;
                  active_thread[(617*4)+3] <= 1'b1;
                  spc617_inst_done         <= `ARIANE_CORE617.piton_pc_vld;
                  spc617_phy_pc_w          <= `ARIANE_CORE617.piton_pc;
                end
            end
    

            assign spc618_thread_id = 2'b00;
            assign spc618_rtl_pc = spc618_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(618*4)]   <= 1'b0;
                  active_thread[(618*4)+1] <= 1'b0;
                  active_thread[(618*4)+2] <= 1'b0;
                  active_thread[(618*4)+3] <= 1'b0;
                  spc618_inst_done         <= 0;
                  spc618_phy_pc_w          <= 0;
                end else begin
                  active_thread[(618*4)]   <= 1'b1;
                  active_thread[(618*4)+1] <= 1'b1;
                  active_thread[(618*4)+2] <= 1'b1;
                  active_thread[(618*4)+3] <= 1'b1;
                  spc618_inst_done         <= `ARIANE_CORE618.piton_pc_vld;
                  spc618_phy_pc_w          <= `ARIANE_CORE618.piton_pc;
                end
            end
    

            assign spc619_thread_id = 2'b00;
            assign spc619_rtl_pc = spc619_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(619*4)]   <= 1'b0;
                  active_thread[(619*4)+1] <= 1'b0;
                  active_thread[(619*4)+2] <= 1'b0;
                  active_thread[(619*4)+3] <= 1'b0;
                  spc619_inst_done         <= 0;
                  spc619_phy_pc_w          <= 0;
                end else begin
                  active_thread[(619*4)]   <= 1'b1;
                  active_thread[(619*4)+1] <= 1'b1;
                  active_thread[(619*4)+2] <= 1'b1;
                  active_thread[(619*4)+3] <= 1'b1;
                  spc619_inst_done         <= `ARIANE_CORE619.piton_pc_vld;
                  spc619_phy_pc_w          <= `ARIANE_CORE619.piton_pc;
                end
            end
    

            assign spc620_thread_id = 2'b00;
            assign spc620_rtl_pc = spc620_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(620*4)]   <= 1'b0;
                  active_thread[(620*4)+1] <= 1'b0;
                  active_thread[(620*4)+2] <= 1'b0;
                  active_thread[(620*4)+3] <= 1'b0;
                  spc620_inst_done         <= 0;
                  spc620_phy_pc_w          <= 0;
                end else begin
                  active_thread[(620*4)]   <= 1'b1;
                  active_thread[(620*4)+1] <= 1'b1;
                  active_thread[(620*4)+2] <= 1'b1;
                  active_thread[(620*4)+3] <= 1'b1;
                  spc620_inst_done         <= `ARIANE_CORE620.piton_pc_vld;
                  spc620_phy_pc_w          <= `ARIANE_CORE620.piton_pc;
                end
            end
    

            assign spc621_thread_id = 2'b00;
            assign spc621_rtl_pc = spc621_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(621*4)]   <= 1'b0;
                  active_thread[(621*4)+1] <= 1'b0;
                  active_thread[(621*4)+2] <= 1'b0;
                  active_thread[(621*4)+3] <= 1'b0;
                  spc621_inst_done         <= 0;
                  spc621_phy_pc_w          <= 0;
                end else begin
                  active_thread[(621*4)]   <= 1'b1;
                  active_thread[(621*4)+1] <= 1'b1;
                  active_thread[(621*4)+2] <= 1'b1;
                  active_thread[(621*4)+3] <= 1'b1;
                  spc621_inst_done         <= `ARIANE_CORE621.piton_pc_vld;
                  spc621_phy_pc_w          <= `ARIANE_CORE621.piton_pc;
                end
            end
    

            assign spc622_thread_id = 2'b00;
            assign spc622_rtl_pc = spc622_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(622*4)]   <= 1'b0;
                  active_thread[(622*4)+1] <= 1'b0;
                  active_thread[(622*4)+2] <= 1'b0;
                  active_thread[(622*4)+3] <= 1'b0;
                  spc622_inst_done         <= 0;
                  spc622_phy_pc_w          <= 0;
                end else begin
                  active_thread[(622*4)]   <= 1'b1;
                  active_thread[(622*4)+1] <= 1'b1;
                  active_thread[(622*4)+2] <= 1'b1;
                  active_thread[(622*4)+3] <= 1'b1;
                  spc622_inst_done         <= `ARIANE_CORE622.piton_pc_vld;
                  spc622_phy_pc_w          <= `ARIANE_CORE622.piton_pc;
                end
            end
    

            assign spc623_thread_id = 2'b00;
            assign spc623_rtl_pc = spc623_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(623*4)]   <= 1'b0;
                  active_thread[(623*4)+1] <= 1'b0;
                  active_thread[(623*4)+2] <= 1'b0;
                  active_thread[(623*4)+3] <= 1'b0;
                  spc623_inst_done         <= 0;
                  spc623_phy_pc_w          <= 0;
                end else begin
                  active_thread[(623*4)]   <= 1'b1;
                  active_thread[(623*4)+1] <= 1'b1;
                  active_thread[(623*4)+2] <= 1'b1;
                  active_thread[(623*4)+3] <= 1'b1;
                  spc623_inst_done         <= `ARIANE_CORE623.piton_pc_vld;
                  spc623_phy_pc_w          <= `ARIANE_CORE623.piton_pc;
                end
            end
    

            assign spc624_thread_id = 2'b00;
            assign spc624_rtl_pc = spc624_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(624*4)]   <= 1'b0;
                  active_thread[(624*4)+1] <= 1'b0;
                  active_thread[(624*4)+2] <= 1'b0;
                  active_thread[(624*4)+3] <= 1'b0;
                  spc624_inst_done         <= 0;
                  spc624_phy_pc_w          <= 0;
                end else begin
                  active_thread[(624*4)]   <= 1'b1;
                  active_thread[(624*4)+1] <= 1'b1;
                  active_thread[(624*4)+2] <= 1'b1;
                  active_thread[(624*4)+3] <= 1'b1;
                  spc624_inst_done         <= `ARIANE_CORE624.piton_pc_vld;
                  spc624_phy_pc_w          <= `ARIANE_CORE624.piton_pc;
                end
            end
    

            assign spc625_thread_id = 2'b00;
            assign spc625_rtl_pc = spc625_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(625*4)]   <= 1'b0;
                  active_thread[(625*4)+1] <= 1'b0;
                  active_thread[(625*4)+2] <= 1'b0;
                  active_thread[(625*4)+3] <= 1'b0;
                  spc625_inst_done         <= 0;
                  spc625_phy_pc_w          <= 0;
                end else begin
                  active_thread[(625*4)]   <= 1'b1;
                  active_thread[(625*4)+1] <= 1'b1;
                  active_thread[(625*4)+2] <= 1'b1;
                  active_thread[(625*4)+3] <= 1'b1;
                  spc625_inst_done         <= `ARIANE_CORE625.piton_pc_vld;
                  spc625_phy_pc_w          <= `ARIANE_CORE625.piton_pc;
                end
            end
    

            assign spc626_thread_id = 2'b00;
            assign spc626_rtl_pc = spc626_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(626*4)]   <= 1'b0;
                  active_thread[(626*4)+1] <= 1'b0;
                  active_thread[(626*4)+2] <= 1'b0;
                  active_thread[(626*4)+3] <= 1'b0;
                  spc626_inst_done         <= 0;
                  spc626_phy_pc_w          <= 0;
                end else begin
                  active_thread[(626*4)]   <= 1'b1;
                  active_thread[(626*4)+1] <= 1'b1;
                  active_thread[(626*4)+2] <= 1'b1;
                  active_thread[(626*4)+3] <= 1'b1;
                  spc626_inst_done         <= `ARIANE_CORE626.piton_pc_vld;
                  spc626_phy_pc_w          <= `ARIANE_CORE626.piton_pc;
                end
            end
    

            assign spc627_thread_id = 2'b00;
            assign spc627_rtl_pc = spc627_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(627*4)]   <= 1'b0;
                  active_thread[(627*4)+1] <= 1'b0;
                  active_thread[(627*4)+2] <= 1'b0;
                  active_thread[(627*4)+3] <= 1'b0;
                  spc627_inst_done         <= 0;
                  spc627_phy_pc_w          <= 0;
                end else begin
                  active_thread[(627*4)]   <= 1'b1;
                  active_thread[(627*4)+1] <= 1'b1;
                  active_thread[(627*4)+2] <= 1'b1;
                  active_thread[(627*4)+3] <= 1'b1;
                  spc627_inst_done         <= `ARIANE_CORE627.piton_pc_vld;
                  spc627_phy_pc_w          <= `ARIANE_CORE627.piton_pc;
                end
            end
    

            assign spc628_thread_id = 2'b00;
            assign spc628_rtl_pc = spc628_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(628*4)]   <= 1'b0;
                  active_thread[(628*4)+1] <= 1'b0;
                  active_thread[(628*4)+2] <= 1'b0;
                  active_thread[(628*4)+3] <= 1'b0;
                  spc628_inst_done         <= 0;
                  spc628_phy_pc_w          <= 0;
                end else begin
                  active_thread[(628*4)]   <= 1'b1;
                  active_thread[(628*4)+1] <= 1'b1;
                  active_thread[(628*4)+2] <= 1'b1;
                  active_thread[(628*4)+3] <= 1'b1;
                  spc628_inst_done         <= `ARIANE_CORE628.piton_pc_vld;
                  spc628_phy_pc_w          <= `ARIANE_CORE628.piton_pc;
                end
            end
    

            assign spc629_thread_id = 2'b00;
            assign spc629_rtl_pc = spc629_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(629*4)]   <= 1'b0;
                  active_thread[(629*4)+1] <= 1'b0;
                  active_thread[(629*4)+2] <= 1'b0;
                  active_thread[(629*4)+3] <= 1'b0;
                  spc629_inst_done         <= 0;
                  spc629_phy_pc_w          <= 0;
                end else begin
                  active_thread[(629*4)]   <= 1'b1;
                  active_thread[(629*4)+1] <= 1'b1;
                  active_thread[(629*4)+2] <= 1'b1;
                  active_thread[(629*4)+3] <= 1'b1;
                  spc629_inst_done         <= `ARIANE_CORE629.piton_pc_vld;
                  spc629_phy_pc_w          <= `ARIANE_CORE629.piton_pc;
                end
            end
    

            assign spc630_thread_id = 2'b00;
            assign spc630_rtl_pc = spc630_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(630*4)]   <= 1'b0;
                  active_thread[(630*4)+1] <= 1'b0;
                  active_thread[(630*4)+2] <= 1'b0;
                  active_thread[(630*4)+3] <= 1'b0;
                  spc630_inst_done         <= 0;
                  spc630_phy_pc_w          <= 0;
                end else begin
                  active_thread[(630*4)]   <= 1'b1;
                  active_thread[(630*4)+1] <= 1'b1;
                  active_thread[(630*4)+2] <= 1'b1;
                  active_thread[(630*4)+3] <= 1'b1;
                  spc630_inst_done         <= `ARIANE_CORE630.piton_pc_vld;
                  spc630_phy_pc_w          <= `ARIANE_CORE630.piton_pc;
                end
            end
    

            assign spc631_thread_id = 2'b00;
            assign spc631_rtl_pc = spc631_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(631*4)]   <= 1'b0;
                  active_thread[(631*4)+1] <= 1'b0;
                  active_thread[(631*4)+2] <= 1'b0;
                  active_thread[(631*4)+3] <= 1'b0;
                  spc631_inst_done         <= 0;
                  spc631_phy_pc_w          <= 0;
                end else begin
                  active_thread[(631*4)]   <= 1'b1;
                  active_thread[(631*4)+1] <= 1'b1;
                  active_thread[(631*4)+2] <= 1'b1;
                  active_thread[(631*4)+3] <= 1'b1;
                  spc631_inst_done         <= `ARIANE_CORE631.piton_pc_vld;
                  spc631_phy_pc_w          <= `ARIANE_CORE631.piton_pc;
                end
            end
    

            assign spc632_thread_id = 2'b00;
            assign spc632_rtl_pc = spc632_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(632*4)]   <= 1'b0;
                  active_thread[(632*4)+1] <= 1'b0;
                  active_thread[(632*4)+2] <= 1'b0;
                  active_thread[(632*4)+3] <= 1'b0;
                  spc632_inst_done         <= 0;
                  spc632_phy_pc_w          <= 0;
                end else begin
                  active_thread[(632*4)]   <= 1'b1;
                  active_thread[(632*4)+1] <= 1'b1;
                  active_thread[(632*4)+2] <= 1'b1;
                  active_thread[(632*4)+3] <= 1'b1;
                  spc632_inst_done         <= `ARIANE_CORE632.piton_pc_vld;
                  spc632_phy_pc_w          <= `ARIANE_CORE632.piton_pc;
                end
            end
    

            assign spc633_thread_id = 2'b00;
            assign spc633_rtl_pc = spc633_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(633*4)]   <= 1'b0;
                  active_thread[(633*4)+1] <= 1'b0;
                  active_thread[(633*4)+2] <= 1'b0;
                  active_thread[(633*4)+3] <= 1'b0;
                  spc633_inst_done         <= 0;
                  spc633_phy_pc_w          <= 0;
                end else begin
                  active_thread[(633*4)]   <= 1'b1;
                  active_thread[(633*4)+1] <= 1'b1;
                  active_thread[(633*4)+2] <= 1'b1;
                  active_thread[(633*4)+3] <= 1'b1;
                  spc633_inst_done         <= `ARIANE_CORE633.piton_pc_vld;
                  spc633_phy_pc_w          <= `ARIANE_CORE633.piton_pc;
                end
            end
    

            assign spc634_thread_id = 2'b00;
            assign spc634_rtl_pc = spc634_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(634*4)]   <= 1'b0;
                  active_thread[(634*4)+1] <= 1'b0;
                  active_thread[(634*4)+2] <= 1'b0;
                  active_thread[(634*4)+3] <= 1'b0;
                  spc634_inst_done         <= 0;
                  spc634_phy_pc_w          <= 0;
                end else begin
                  active_thread[(634*4)]   <= 1'b1;
                  active_thread[(634*4)+1] <= 1'b1;
                  active_thread[(634*4)+2] <= 1'b1;
                  active_thread[(634*4)+3] <= 1'b1;
                  spc634_inst_done         <= `ARIANE_CORE634.piton_pc_vld;
                  spc634_phy_pc_w          <= `ARIANE_CORE634.piton_pc;
                end
            end
    

            assign spc635_thread_id = 2'b00;
            assign spc635_rtl_pc = spc635_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(635*4)]   <= 1'b0;
                  active_thread[(635*4)+1] <= 1'b0;
                  active_thread[(635*4)+2] <= 1'b0;
                  active_thread[(635*4)+3] <= 1'b0;
                  spc635_inst_done         <= 0;
                  spc635_phy_pc_w          <= 0;
                end else begin
                  active_thread[(635*4)]   <= 1'b1;
                  active_thread[(635*4)+1] <= 1'b1;
                  active_thread[(635*4)+2] <= 1'b1;
                  active_thread[(635*4)+3] <= 1'b1;
                  spc635_inst_done         <= `ARIANE_CORE635.piton_pc_vld;
                  spc635_phy_pc_w          <= `ARIANE_CORE635.piton_pc;
                end
            end
    

            assign spc636_thread_id = 2'b00;
            assign spc636_rtl_pc = spc636_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(636*4)]   <= 1'b0;
                  active_thread[(636*4)+1] <= 1'b0;
                  active_thread[(636*4)+2] <= 1'b0;
                  active_thread[(636*4)+3] <= 1'b0;
                  spc636_inst_done         <= 0;
                  spc636_phy_pc_w          <= 0;
                end else begin
                  active_thread[(636*4)]   <= 1'b1;
                  active_thread[(636*4)+1] <= 1'b1;
                  active_thread[(636*4)+2] <= 1'b1;
                  active_thread[(636*4)+3] <= 1'b1;
                  spc636_inst_done         <= `ARIANE_CORE636.piton_pc_vld;
                  spc636_phy_pc_w          <= `ARIANE_CORE636.piton_pc;
                end
            end
    

            assign spc637_thread_id = 2'b00;
            assign spc637_rtl_pc = spc637_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(637*4)]   <= 1'b0;
                  active_thread[(637*4)+1] <= 1'b0;
                  active_thread[(637*4)+2] <= 1'b0;
                  active_thread[(637*4)+3] <= 1'b0;
                  spc637_inst_done         <= 0;
                  spc637_phy_pc_w          <= 0;
                end else begin
                  active_thread[(637*4)]   <= 1'b1;
                  active_thread[(637*4)+1] <= 1'b1;
                  active_thread[(637*4)+2] <= 1'b1;
                  active_thread[(637*4)+3] <= 1'b1;
                  spc637_inst_done         <= `ARIANE_CORE637.piton_pc_vld;
                  spc637_phy_pc_w          <= `ARIANE_CORE637.piton_pc;
                end
            end
    

            assign spc638_thread_id = 2'b00;
            assign spc638_rtl_pc = spc638_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(638*4)]   <= 1'b0;
                  active_thread[(638*4)+1] <= 1'b0;
                  active_thread[(638*4)+2] <= 1'b0;
                  active_thread[(638*4)+3] <= 1'b0;
                  spc638_inst_done         <= 0;
                  spc638_phy_pc_w          <= 0;
                end else begin
                  active_thread[(638*4)]   <= 1'b1;
                  active_thread[(638*4)+1] <= 1'b1;
                  active_thread[(638*4)+2] <= 1'b1;
                  active_thread[(638*4)+3] <= 1'b1;
                  spc638_inst_done         <= `ARIANE_CORE638.piton_pc_vld;
                  spc638_phy_pc_w          <= `ARIANE_CORE638.piton_pc;
                end
            end
    

            assign spc639_thread_id = 2'b00;
            assign spc639_rtl_pc = spc639_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(639*4)]   <= 1'b0;
                  active_thread[(639*4)+1] <= 1'b0;
                  active_thread[(639*4)+2] <= 1'b0;
                  active_thread[(639*4)+3] <= 1'b0;
                  spc639_inst_done         <= 0;
                  spc639_phy_pc_w          <= 0;
                end else begin
                  active_thread[(639*4)]   <= 1'b1;
                  active_thread[(639*4)+1] <= 1'b1;
                  active_thread[(639*4)+2] <= 1'b1;
                  active_thread[(639*4)+3] <= 1'b1;
                  spc639_inst_done         <= `ARIANE_CORE639.piton_pc_vld;
                  spc639_phy_pc_w          <= `ARIANE_CORE639.piton_pc;
                end
            end
    

            assign spc640_thread_id = 2'b00;
            assign spc640_rtl_pc = spc640_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(640*4)]   <= 1'b0;
                  active_thread[(640*4)+1] <= 1'b0;
                  active_thread[(640*4)+2] <= 1'b0;
                  active_thread[(640*4)+3] <= 1'b0;
                  spc640_inst_done         <= 0;
                  spc640_phy_pc_w          <= 0;
                end else begin
                  active_thread[(640*4)]   <= 1'b1;
                  active_thread[(640*4)+1] <= 1'b1;
                  active_thread[(640*4)+2] <= 1'b1;
                  active_thread[(640*4)+3] <= 1'b1;
                  spc640_inst_done         <= `ARIANE_CORE640.piton_pc_vld;
                  spc640_phy_pc_w          <= `ARIANE_CORE640.piton_pc;
                end
            end
    

            assign spc641_thread_id = 2'b00;
            assign spc641_rtl_pc = spc641_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(641*4)]   <= 1'b0;
                  active_thread[(641*4)+1] <= 1'b0;
                  active_thread[(641*4)+2] <= 1'b0;
                  active_thread[(641*4)+3] <= 1'b0;
                  spc641_inst_done         <= 0;
                  spc641_phy_pc_w          <= 0;
                end else begin
                  active_thread[(641*4)]   <= 1'b1;
                  active_thread[(641*4)+1] <= 1'b1;
                  active_thread[(641*4)+2] <= 1'b1;
                  active_thread[(641*4)+3] <= 1'b1;
                  spc641_inst_done         <= `ARIANE_CORE641.piton_pc_vld;
                  spc641_phy_pc_w          <= `ARIANE_CORE641.piton_pc;
                end
            end
    

            assign spc642_thread_id = 2'b00;
            assign spc642_rtl_pc = spc642_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(642*4)]   <= 1'b0;
                  active_thread[(642*4)+1] <= 1'b0;
                  active_thread[(642*4)+2] <= 1'b0;
                  active_thread[(642*4)+3] <= 1'b0;
                  spc642_inst_done         <= 0;
                  spc642_phy_pc_w          <= 0;
                end else begin
                  active_thread[(642*4)]   <= 1'b1;
                  active_thread[(642*4)+1] <= 1'b1;
                  active_thread[(642*4)+2] <= 1'b1;
                  active_thread[(642*4)+3] <= 1'b1;
                  spc642_inst_done         <= `ARIANE_CORE642.piton_pc_vld;
                  spc642_phy_pc_w          <= `ARIANE_CORE642.piton_pc;
                end
            end
    

            assign spc643_thread_id = 2'b00;
            assign spc643_rtl_pc = spc643_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(643*4)]   <= 1'b0;
                  active_thread[(643*4)+1] <= 1'b0;
                  active_thread[(643*4)+2] <= 1'b0;
                  active_thread[(643*4)+3] <= 1'b0;
                  spc643_inst_done         <= 0;
                  spc643_phy_pc_w          <= 0;
                end else begin
                  active_thread[(643*4)]   <= 1'b1;
                  active_thread[(643*4)+1] <= 1'b1;
                  active_thread[(643*4)+2] <= 1'b1;
                  active_thread[(643*4)+3] <= 1'b1;
                  spc643_inst_done         <= `ARIANE_CORE643.piton_pc_vld;
                  spc643_phy_pc_w          <= `ARIANE_CORE643.piton_pc;
                end
            end
    

            assign spc644_thread_id = 2'b00;
            assign spc644_rtl_pc = spc644_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(644*4)]   <= 1'b0;
                  active_thread[(644*4)+1] <= 1'b0;
                  active_thread[(644*4)+2] <= 1'b0;
                  active_thread[(644*4)+3] <= 1'b0;
                  spc644_inst_done         <= 0;
                  spc644_phy_pc_w          <= 0;
                end else begin
                  active_thread[(644*4)]   <= 1'b1;
                  active_thread[(644*4)+1] <= 1'b1;
                  active_thread[(644*4)+2] <= 1'b1;
                  active_thread[(644*4)+3] <= 1'b1;
                  spc644_inst_done         <= `ARIANE_CORE644.piton_pc_vld;
                  spc644_phy_pc_w          <= `ARIANE_CORE644.piton_pc;
                end
            end
    

            assign spc645_thread_id = 2'b00;
            assign spc645_rtl_pc = spc645_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(645*4)]   <= 1'b0;
                  active_thread[(645*4)+1] <= 1'b0;
                  active_thread[(645*4)+2] <= 1'b0;
                  active_thread[(645*4)+3] <= 1'b0;
                  spc645_inst_done         <= 0;
                  spc645_phy_pc_w          <= 0;
                end else begin
                  active_thread[(645*4)]   <= 1'b1;
                  active_thread[(645*4)+1] <= 1'b1;
                  active_thread[(645*4)+2] <= 1'b1;
                  active_thread[(645*4)+3] <= 1'b1;
                  spc645_inst_done         <= `ARIANE_CORE645.piton_pc_vld;
                  spc645_phy_pc_w          <= `ARIANE_CORE645.piton_pc;
                end
            end
    

            assign spc646_thread_id = 2'b00;
            assign spc646_rtl_pc = spc646_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(646*4)]   <= 1'b0;
                  active_thread[(646*4)+1] <= 1'b0;
                  active_thread[(646*4)+2] <= 1'b0;
                  active_thread[(646*4)+3] <= 1'b0;
                  spc646_inst_done         <= 0;
                  spc646_phy_pc_w          <= 0;
                end else begin
                  active_thread[(646*4)]   <= 1'b1;
                  active_thread[(646*4)+1] <= 1'b1;
                  active_thread[(646*4)+2] <= 1'b1;
                  active_thread[(646*4)+3] <= 1'b1;
                  spc646_inst_done         <= `ARIANE_CORE646.piton_pc_vld;
                  spc646_phy_pc_w          <= `ARIANE_CORE646.piton_pc;
                end
            end
    

            assign spc647_thread_id = 2'b00;
            assign spc647_rtl_pc = spc647_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(647*4)]   <= 1'b0;
                  active_thread[(647*4)+1] <= 1'b0;
                  active_thread[(647*4)+2] <= 1'b0;
                  active_thread[(647*4)+3] <= 1'b0;
                  spc647_inst_done         <= 0;
                  spc647_phy_pc_w          <= 0;
                end else begin
                  active_thread[(647*4)]   <= 1'b1;
                  active_thread[(647*4)+1] <= 1'b1;
                  active_thread[(647*4)+2] <= 1'b1;
                  active_thread[(647*4)+3] <= 1'b1;
                  spc647_inst_done         <= `ARIANE_CORE647.piton_pc_vld;
                  spc647_phy_pc_w          <= `ARIANE_CORE647.piton_pc;
                end
            end
    

            assign spc648_thread_id = 2'b00;
            assign spc648_rtl_pc = spc648_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(648*4)]   <= 1'b0;
                  active_thread[(648*4)+1] <= 1'b0;
                  active_thread[(648*4)+2] <= 1'b0;
                  active_thread[(648*4)+3] <= 1'b0;
                  spc648_inst_done         <= 0;
                  spc648_phy_pc_w          <= 0;
                end else begin
                  active_thread[(648*4)]   <= 1'b1;
                  active_thread[(648*4)+1] <= 1'b1;
                  active_thread[(648*4)+2] <= 1'b1;
                  active_thread[(648*4)+3] <= 1'b1;
                  spc648_inst_done         <= `ARIANE_CORE648.piton_pc_vld;
                  spc648_phy_pc_w          <= `ARIANE_CORE648.piton_pc;
                end
            end
    

            assign spc649_thread_id = 2'b00;
            assign spc649_rtl_pc = spc649_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(649*4)]   <= 1'b0;
                  active_thread[(649*4)+1] <= 1'b0;
                  active_thread[(649*4)+2] <= 1'b0;
                  active_thread[(649*4)+3] <= 1'b0;
                  spc649_inst_done         <= 0;
                  spc649_phy_pc_w          <= 0;
                end else begin
                  active_thread[(649*4)]   <= 1'b1;
                  active_thread[(649*4)+1] <= 1'b1;
                  active_thread[(649*4)+2] <= 1'b1;
                  active_thread[(649*4)+3] <= 1'b1;
                  spc649_inst_done         <= `ARIANE_CORE649.piton_pc_vld;
                  spc649_phy_pc_w          <= `ARIANE_CORE649.piton_pc;
                end
            end
    

            assign spc650_thread_id = 2'b00;
            assign spc650_rtl_pc = spc650_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(650*4)]   <= 1'b0;
                  active_thread[(650*4)+1] <= 1'b0;
                  active_thread[(650*4)+2] <= 1'b0;
                  active_thread[(650*4)+3] <= 1'b0;
                  spc650_inst_done         <= 0;
                  spc650_phy_pc_w          <= 0;
                end else begin
                  active_thread[(650*4)]   <= 1'b1;
                  active_thread[(650*4)+1] <= 1'b1;
                  active_thread[(650*4)+2] <= 1'b1;
                  active_thread[(650*4)+3] <= 1'b1;
                  spc650_inst_done         <= `ARIANE_CORE650.piton_pc_vld;
                  spc650_phy_pc_w          <= `ARIANE_CORE650.piton_pc;
                end
            end
    

            assign spc651_thread_id = 2'b00;
            assign spc651_rtl_pc = spc651_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(651*4)]   <= 1'b0;
                  active_thread[(651*4)+1] <= 1'b0;
                  active_thread[(651*4)+2] <= 1'b0;
                  active_thread[(651*4)+3] <= 1'b0;
                  spc651_inst_done         <= 0;
                  spc651_phy_pc_w          <= 0;
                end else begin
                  active_thread[(651*4)]   <= 1'b1;
                  active_thread[(651*4)+1] <= 1'b1;
                  active_thread[(651*4)+2] <= 1'b1;
                  active_thread[(651*4)+3] <= 1'b1;
                  spc651_inst_done         <= `ARIANE_CORE651.piton_pc_vld;
                  spc651_phy_pc_w          <= `ARIANE_CORE651.piton_pc;
                end
            end
    

            assign spc652_thread_id = 2'b00;
            assign spc652_rtl_pc = spc652_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(652*4)]   <= 1'b0;
                  active_thread[(652*4)+1] <= 1'b0;
                  active_thread[(652*4)+2] <= 1'b0;
                  active_thread[(652*4)+3] <= 1'b0;
                  spc652_inst_done         <= 0;
                  spc652_phy_pc_w          <= 0;
                end else begin
                  active_thread[(652*4)]   <= 1'b1;
                  active_thread[(652*4)+1] <= 1'b1;
                  active_thread[(652*4)+2] <= 1'b1;
                  active_thread[(652*4)+3] <= 1'b1;
                  spc652_inst_done         <= `ARIANE_CORE652.piton_pc_vld;
                  spc652_phy_pc_w          <= `ARIANE_CORE652.piton_pc;
                end
            end
    

            assign spc653_thread_id = 2'b00;
            assign spc653_rtl_pc = spc653_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(653*4)]   <= 1'b0;
                  active_thread[(653*4)+1] <= 1'b0;
                  active_thread[(653*4)+2] <= 1'b0;
                  active_thread[(653*4)+3] <= 1'b0;
                  spc653_inst_done         <= 0;
                  spc653_phy_pc_w          <= 0;
                end else begin
                  active_thread[(653*4)]   <= 1'b1;
                  active_thread[(653*4)+1] <= 1'b1;
                  active_thread[(653*4)+2] <= 1'b1;
                  active_thread[(653*4)+3] <= 1'b1;
                  spc653_inst_done         <= `ARIANE_CORE653.piton_pc_vld;
                  spc653_phy_pc_w          <= `ARIANE_CORE653.piton_pc;
                end
            end
    

            assign spc654_thread_id = 2'b00;
            assign spc654_rtl_pc = spc654_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(654*4)]   <= 1'b0;
                  active_thread[(654*4)+1] <= 1'b0;
                  active_thread[(654*4)+2] <= 1'b0;
                  active_thread[(654*4)+3] <= 1'b0;
                  spc654_inst_done         <= 0;
                  spc654_phy_pc_w          <= 0;
                end else begin
                  active_thread[(654*4)]   <= 1'b1;
                  active_thread[(654*4)+1] <= 1'b1;
                  active_thread[(654*4)+2] <= 1'b1;
                  active_thread[(654*4)+3] <= 1'b1;
                  spc654_inst_done         <= `ARIANE_CORE654.piton_pc_vld;
                  spc654_phy_pc_w          <= `ARIANE_CORE654.piton_pc;
                end
            end
    

            assign spc655_thread_id = 2'b00;
            assign spc655_rtl_pc = spc655_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(655*4)]   <= 1'b0;
                  active_thread[(655*4)+1] <= 1'b0;
                  active_thread[(655*4)+2] <= 1'b0;
                  active_thread[(655*4)+3] <= 1'b0;
                  spc655_inst_done         <= 0;
                  spc655_phy_pc_w          <= 0;
                end else begin
                  active_thread[(655*4)]   <= 1'b1;
                  active_thread[(655*4)+1] <= 1'b1;
                  active_thread[(655*4)+2] <= 1'b1;
                  active_thread[(655*4)+3] <= 1'b1;
                  spc655_inst_done         <= `ARIANE_CORE655.piton_pc_vld;
                  spc655_phy_pc_w          <= `ARIANE_CORE655.piton_pc;
                end
            end
    

            assign spc656_thread_id = 2'b00;
            assign spc656_rtl_pc = spc656_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(656*4)]   <= 1'b0;
                  active_thread[(656*4)+1] <= 1'b0;
                  active_thread[(656*4)+2] <= 1'b0;
                  active_thread[(656*4)+3] <= 1'b0;
                  spc656_inst_done         <= 0;
                  spc656_phy_pc_w          <= 0;
                end else begin
                  active_thread[(656*4)]   <= 1'b1;
                  active_thread[(656*4)+1] <= 1'b1;
                  active_thread[(656*4)+2] <= 1'b1;
                  active_thread[(656*4)+3] <= 1'b1;
                  spc656_inst_done         <= `ARIANE_CORE656.piton_pc_vld;
                  spc656_phy_pc_w          <= `ARIANE_CORE656.piton_pc;
                end
            end
    

            assign spc657_thread_id = 2'b00;
            assign spc657_rtl_pc = spc657_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(657*4)]   <= 1'b0;
                  active_thread[(657*4)+1] <= 1'b0;
                  active_thread[(657*4)+2] <= 1'b0;
                  active_thread[(657*4)+3] <= 1'b0;
                  spc657_inst_done         <= 0;
                  spc657_phy_pc_w          <= 0;
                end else begin
                  active_thread[(657*4)]   <= 1'b1;
                  active_thread[(657*4)+1] <= 1'b1;
                  active_thread[(657*4)+2] <= 1'b1;
                  active_thread[(657*4)+3] <= 1'b1;
                  spc657_inst_done         <= `ARIANE_CORE657.piton_pc_vld;
                  spc657_phy_pc_w          <= `ARIANE_CORE657.piton_pc;
                end
            end
    

            assign spc658_thread_id = 2'b00;
            assign spc658_rtl_pc = spc658_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(658*4)]   <= 1'b0;
                  active_thread[(658*4)+1] <= 1'b0;
                  active_thread[(658*4)+2] <= 1'b0;
                  active_thread[(658*4)+3] <= 1'b0;
                  spc658_inst_done         <= 0;
                  spc658_phy_pc_w          <= 0;
                end else begin
                  active_thread[(658*4)]   <= 1'b1;
                  active_thread[(658*4)+1] <= 1'b1;
                  active_thread[(658*4)+2] <= 1'b1;
                  active_thread[(658*4)+3] <= 1'b1;
                  spc658_inst_done         <= `ARIANE_CORE658.piton_pc_vld;
                  spc658_phy_pc_w          <= `ARIANE_CORE658.piton_pc;
                end
            end
    

            assign spc659_thread_id = 2'b00;
            assign spc659_rtl_pc = spc659_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(659*4)]   <= 1'b0;
                  active_thread[(659*4)+1] <= 1'b0;
                  active_thread[(659*4)+2] <= 1'b0;
                  active_thread[(659*4)+3] <= 1'b0;
                  spc659_inst_done         <= 0;
                  spc659_phy_pc_w          <= 0;
                end else begin
                  active_thread[(659*4)]   <= 1'b1;
                  active_thread[(659*4)+1] <= 1'b1;
                  active_thread[(659*4)+2] <= 1'b1;
                  active_thread[(659*4)+3] <= 1'b1;
                  spc659_inst_done         <= `ARIANE_CORE659.piton_pc_vld;
                  spc659_phy_pc_w          <= `ARIANE_CORE659.piton_pc;
                end
            end
    

            assign spc660_thread_id = 2'b00;
            assign spc660_rtl_pc = spc660_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(660*4)]   <= 1'b0;
                  active_thread[(660*4)+1] <= 1'b0;
                  active_thread[(660*4)+2] <= 1'b0;
                  active_thread[(660*4)+3] <= 1'b0;
                  spc660_inst_done         <= 0;
                  spc660_phy_pc_w          <= 0;
                end else begin
                  active_thread[(660*4)]   <= 1'b1;
                  active_thread[(660*4)+1] <= 1'b1;
                  active_thread[(660*4)+2] <= 1'b1;
                  active_thread[(660*4)+3] <= 1'b1;
                  spc660_inst_done         <= `ARIANE_CORE660.piton_pc_vld;
                  spc660_phy_pc_w          <= `ARIANE_CORE660.piton_pc;
                end
            end
    

            assign spc661_thread_id = 2'b00;
            assign spc661_rtl_pc = spc661_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(661*4)]   <= 1'b0;
                  active_thread[(661*4)+1] <= 1'b0;
                  active_thread[(661*4)+2] <= 1'b0;
                  active_thread[(661*4)+3] <= 1'b0;
                  spc661_inst_done         <= 0;
                  spc661_phy_pc_w          <= 0;
                end else begin
                  active_thread[(661*4)]   <= 1'b1;
                  active_thread[(661*4)+1] <= 1'b1;
                  active_thread[(661*4)+2] <= 1'b1;
                  active_thread[(661*4)+3] <= 1'b1;
                  spc661_inst_done         <= `ARIANE_CORE661.piton_pc_vld;
                  spc661_phy_pc_w          <= `ARIANE_CORE661.piton_pc;
                end
            end
    

            assign spc662_thread_id = 2'b00;
            assign spc662_rtl_pc = spc662_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(662*4)]   <= 1'b0;
                  active_thread[(662*4)+1] <= 1'b0;
                  active_thread[(662*4)+2] <= 1'b0;
                  active_thread[(662*4)+3] <= 1'b0;
                  spc662_inst_done         <= 0;
                  spc662_phy_pc_w          <= 0;
                end else begin
                  active_thread[(662*4)]   <= 1'b1;
                  active_thread[(662*4)+1] <= 1'b1;
                  active_thread[(662*4)+2] <= 1'b1;
                  active_thread[(662*4)+3] <= 1'b1;
                  spc662_inst_done         <= `ARIANE_CORE662.piton_pc_vld;
                  spc662_phy_pc_w          <= `ARIANE_CORE662.piton_pc;
                end
            end
    

            assign spc663_thread_id = 2'b00;
            assign spc663_rtl_pc = spc663_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(663*4)]   <= 1'b0;
                  active_thread[(663*4)+1] <= 1'b0;
                  active_thread[(663*4)+2] <= 1'b0;
                  active_thread[(663*4)+3] <= 1'b0;
                  spc663_inst_done         <= 0;
                  spc663_phy_pc_w          <= 0;
                end else begin
                  active_thread[(663*4)]   <= 1'b1;
                  active_thread[(663*4)+1] <= 1'b1;
                  active_thread[(663*4)+2] <= 1'b1;
                  active_thread[(663*4)+3] <= 1'b1;
                  spc663_inst_done         <= `ARIANE_CORE663.piton_pc_vld;
                  spc663_phy_pc_w          <= `ARIANE_CORE663.piton_pc;
                end
            end
    

            assign spc664_thread_id = 2'b00;
            assign spc664_rtl_pc = spc664_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(664*4)]   <= 1'b0;
                  active_thread[(664*4)+1] <= 1'b0;
                  active_thread[(664*4)+2] <= 1'b0;
                  active_thread[(664*4)+3] <= 1'b0;
                  spc664_inst_done         <= 0;
                  spc664_phy_pc_w          <= 0;
                end else begin
                  active_thread[(664*4)]   <= 1'b1;
                  active_thread[(664*4)+1] <= 1'b1;
                  active_thread[(664*4)+2] <= 1'b1;
                  active_thread[(664*4)+3] <= 1'b1;
                  spc664_inst_done         <= `ARIANE_CORE664.piton_pc_vld;
                  spc664_phy_pc_w          <= `ARIANE_CORE664.piton_pc;
                end
            end
    

            assign spc665_thread_id = 2'b00;
            assign spc665_rtl_pc = spc665_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(665*4)]   <= 1'b0;
                  active_thread[(665*4)+1] <= 1'b0;
                  active_thread[(665*4)+2] <= 1'b0;
                  active_thread[(665*4)+3] <= 1'b0;
                  spc665_inst_done         <= 0;
                  spc665_phy_pc_w          <= 0;
                end else begin
                  active_thread[(665*4)]   <= 1'b1;
                  active_thread[(665*4)+1] <= 1'b1;
                  active_thread[(665*4)+2] <= 1'b1;
                  active_thread[(665*4)+3] <= 1'b1;
                  spc665_inst_done         <= `ARIANE_CORE665.piton_pc_vld;
                  spc665_phy_pc_w          <= `ARIANE_CORE665.piton_pc;
                end
            end
    

            assign spc666_thread_id = 2'b00;
            assign spc666_rtl_pc = spc666_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(666*4)]   <= 1'b0;
                  active_thread[(666*4)+1] <= 1'b0;
                  active_thread[(666*4)+2] <= 1'b0;
                  active_thread[(666*4)+3] <= 1'b0;
                  spc666_inst_done         <= 0;
                  spc666_phy_pc_w          <= 0;
                end else begin
                  active_thread[(666*4)]   <= 1'b1;
                  active_thread[(666*4)+1] <= 1'b1;
                  active_thread[(666*4)+2] <= 1'b1;
                  active_thread[(666*4)+3] <= 1'b1;
                  spc666_inst_done         <= `ARIANE_CORE666.piton_pc_vld;
                  spc666_phy_pc_w          <= `ARIANE_CORE666.piton_pc;
                end
            end
    

            assign spc667_thread_id = 2'b00;
            assign spc667_rtl_pc = spc667_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(667*4)]   <= 1'b0;
                  active_thread[(667*4)+1] <= 1'b0;
                  active_thread[(667*4)+2] <= 1'b0;
                  active_thread[(667*4)+3] <= 1'b0;
                  spc667_inst_done         <= 0;
                  spc667_phy_pc_w          <= 0;
                end else begin
                  active_thread[(667*4)]   <= 1'b1;
                  active_thread[(667*4)+1] <= 1'b1;
                  active_thread[(667*4)+2] <= 1'b1;
                  active_thread[(667*4)+3] <= 1'b1;
                  spc667_inst_done         <= `ARIANE_CORE667.piton_pc_vld;
                  spc667_phy_pc_w          <= `ARIANE_CORE667.piton_pc;
                end
            end
    

            assign spc668_thread_id = 2'b00;
            assign spc668_rtl_pc = spc668_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(668*4)]   <= 1'b0;
                  active_thread[(668*4)+1] <= 1'b0;
                  active_thread[(668*4)+2] <= 1'b0;
                  active_thread[(668*4)+3] <= 1'b0;
                  spc668_inst_done         <= 0;
                  spc668_phy_pc_w          <= 0;
                end else begin
                  active_thread[(668*4)]   <= 1'b1;
                  active_thread[(668*4)+1] <= 1'b1;
                  active_thread[(668*4)+2] <= 1'b1;
                  active_thread[(668*4)+3] <= 1'b1;
                  spc668_inst_done         <= `ARIANE_CORE668.piton_pc_vld;
                  spc668_phy_pc_w          <= `ARIANE_CORE668.piton_pc;
                end
            end
    

            assign spc669_thread_id = 2'b00;
            assign spc669_rtl_pc = spc669_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(669*4)]   <= 1'b0;
                  active_thread[(669*4)+1] <= 1'b0;
                  active_thread[(669*4)+2] <= 1'b0;
                  active_thread[(669*4)+3] <= 1'b0;
                  spc669_inst_done         <= 0;
                  spc669_phy_pc_w          <= 0;
                end else begin
                  active_thread[(669*4)]   <= 1'b1;
                  active_thread[(669*4)+1] <= 1'b1;
                  active_thread[(669*4)+2] <= 1'b1;
                  active_thread[(669*4)+3] <= 1'b1;
                  spc669_inst_done         <= `ARIANE_CORE669.piton_pc_vld;
                  spc669_phy_pc_w          <= `ARIANE_CORE669.piton_pc;
                end
            end
    

            assign spc670_thread_id = 2'b00;
            assign spc670_rtl_pc = spc670_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(670*4)]   <= 1'b0;
                  active_thread[(670*4)+1] <= 1'b0;
                  active_thread[(670*4)+2] <= 1'b0;
                  active_thread[(670*4)+3] <= 1'b0;
                  spc670_inst_done         <= 0;
                  spc670_phy_pc_w          <= 0;
                end else begin
                  active_thread[(670*4)]   <= 1'b1;
                  active_thread[(670*4)+1] <= 1'b1;
                  active_thread[(670*4)+2] <= 1'b1;
                  active_thread[(670*4)+3] <= 1'b1;
                  spc670_inst_done         <= `ARIANE_CORE670.piton_pc_vld;
                  spc670_phy_pc_w          <= `ARIANE_CORE670.piton_pc;
                end
            end
    

            assign spc671_thread_id = 2'b00;
            assign spc671_rtl_pc = spc671_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(671*4)]   <= 1'b0;
                  active_thread[(671*4)+1] <= 1'b0;
                  active_thread[(671*4)+2] <= 1'b0;
                  active_thread[(671*4)+3] <= 1'b0;
                  spc671_inst_done         <= 0;
                  spc671_phy_pc_w          <= 0;
                end else begin
                  active_thread[(671*4)]   <= 1'b1;
                  active_thread[(671*4)+1] <= 1'b1;
                  active_thread[(671*4)+2] <= 1'b1;
                  active_thread[(671*4)+3] <= 1'b1;
                  spc671_inst_done         <= `ARIANE_CORE671.piton_pc_vld;
                  spc671_phy_pc_w          <= `ARIANE_CORE671.piton_pc;
                end
            end
    

            assign spc672_thread_id = 2'b00;
            assign spc672_rtl_pc = spc672_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(672*4)]   <= 1'b0;
                  active_thread[(672*4)+1] <= 1'b0;
                  active_thread[(672*4)+2] <= 1'b0;
                  active_thread[(672*4)+3] <= 1'b0;
                  spc672_inst_done         <= 0;
                  spc672_phy_pc_w          <= 0;
                end else begin
                  active_thread[(672*4)]   <= 1'b1;
                  active_thread[(672*4)+1] <= 1'b1;
                  active_thread[(672*4)+2] <= 1'b1;
                  active_thread[(672*4)+3] <= 1'b1;
                  spc672_inst_done         <= `ARIANE_CORE672.piton_pc_vld;
                  spc672_phy_pc_w          <= `ARIANE_CORE672.piton_pc;
                end
            end
    

            assign spc673_thread_id = 2'b00;
            assign spc673_rtl_pc = spc673_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(673*4)]   <= 1'b0;
                  active_thread[(673*4)+1] <= 1'b0;
                  active_thread[(673*4)+2] <= 1'b0;
                  active_thread[(673*4)+3] <= 1'b0;
                  spc673_inst_done         <= 0;
                  spc673_phy_pc_w          <= 0;
                end else begin
                  active_thread[(673*4)]   <= 1'b1;
                  active_thread[(673*4)+1] <= 1'b1;
                  active_thread[(673*4)+2] <= 1'b1;
                  active_thread[(673*4)+3] <= 1'b1;
                  spc673_inst_done         <= `ARIANE_CORE673.piton_pc_vld;
                  spc673_phy_pc_w          <= `ARIANE_CORE673.piton_pc;
                end
            end
    

            assign spc674_thread_id = 2'b00;
            assign spc674_rtl_pc = spc674_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(674*4)]   <= 1'b0;
                  active_thread[(674*4)+1] <= 1'b0;
                  active_thread[(674*4)+2] <= 1'b0;
                  active_thread[(674*4)+3] <= 1'b0;
                  spc674_inst_done         <= 0;
                  spc674_phy_pc_w          <= 0;
                end else begin
                  active_thread[(674*4)]   <= 1'b1;
                  active_thread[(674*4)+1] <= 1'b1;
                  active_thread[(674*4)+2] <= 1'b1;
                  active_thread[(674*4)+3] <= 1'b1;
                  spc674_inst_done         <= `ARIANE_CORE674.piton_pc_vld;
                  spc674_phy_pc_w          <= `ARIANE_CORE674.piton_pc;
                end
            end
    

            assign spc675_thread_id = 2'b00;
            assign spc675_rtl_pc = spc675_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(675*4)]   <= 1'b0;
                  active_thread[(675*4)+1] <= 1'b0;
                  active_thread[(675*4)+2] <= 1'b0;
                  active_thread[(675*4)+3] <= 1'b0;
                  spc675_inst_done         <= 0;
                  spc675_phy_pc_w          <= 0;
                end else begin
                  active_thread[(675*4)]   <= 1'b1;
                  active_thread[(675*4)+1] <= 1'b1;
                  active_thread[(675*4)+2] <= 1'b1;
                  active_thread[(675*4)+3] <= 1'b1;
                  spc675_inst_done         <= `ARIANE_CORE675.piton_pc_vld;
                  spc675_phy_pc_w          <= `ARIANE_CORE675.piton_pc;
                end
            end
    

            assign spc676_thread_id = 2'b00;
            assign spc676_rtl_pc = spc676_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(676*4)]   <= 1'b0;
                  active_thread[(676*4)+1] <= 1'b0;
                  active_thread[(676*4)+2] <= 1'b0;
                  active_thread[(676*4)+3] <= 1'b0;
                  spc676_inst_done         <= 0;
                  spc676_phy_pc_w          <= 0;
                end else begin
                  active_thread[(676*4)]   <= 1'b1;
                  active_thread[(676*4)+1] <= 1'b1;
                  active_thread[(676*4)+2] <= 1'b1;
                  active_thread[(676*4)+3] <= 1'b1;
                  spc676_inst_done         <= `ARIANE_CORE676.piton_pc_vld;
                  spc676_phy_pc_w          <= `ARIANE_CORE676.piton_pc;
                end
            end
    

            assign spc677_thread_id = 2'b00;
            assign spc677_rtl_pc = spc677_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(677*4)]   <= 1'b0;
                  active_thread[(677*4)+1] <= 1'b0;
                  active_thread[(677*4)+2] <= 1'b0;
                  active_thread[(677*4)+3] <= 1'b0;
                  spc677_inst_done         <= 0;
                  spc677_phy_pc_w          <= 0;
                end else begin
                  active_thread[(677*4)]   <= 1'b1;
                  active_thread[(677*4)+1] <= 1'b1;
                  active_thread[(677*4)+2] <= 1'b1;
                  active_thread[(677*4)+3] <= 1'b1;
                  spc677_inst_done         <= `ARIANE_CORE677.piton_pc_vld;
                  spc677_phy_pc_w          <= `ARIANE_CORE677.piton_pc;
                end
            end
    

            assign spc678_thread_id = 2'b00;
            assign spc678_rtl_pc = spc678_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(678*4)]   <= 1'b0;
                  active_thread[(678*4)+1] <= 1'b0;
                  active_thread[(678*4)+2] <= 1'b0;
                  active_thread[(678*4)+3] <= 1'b0;
                  spc678_inst_done         <= 0;
                  spc678_phy_pc_w          <= 0;
                end else begin
                  active_thread[(678*4)]   <= 1'b1;
                  active_thread[(678*4)+1] <= 1'b1;
                  active_thread[(678*4)+2] <= 1'b1;
                  active_thread[(678*4)+3] <= 1'b1;
                  spc678_inst_done         <= `ARIANE_CORE678.piton_pc_vld;
                  spc678_phy_pc_w          <= `ARIANE_CORE678.piton_pc;
                end
            end
    

            assign spc679_thread_id = 2'b00;
            assign spc679_rtl_pc = spc679_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(679*4)]   <= 1'b0;
                  active_thread[(679*4)+1] <= 1'b0;
                  active_thread[(679*4)+2] <= 1'b0;
                  active_thread[(679*4)+3] <= 1'b0;
                  spc679_inst_done         <= 0;
                  spc679_phy_pc_w          <= 0;
                end else begin
                  active_thread[(679*4)]   <= 1'b1;
                  active_thread[(679*4)+1] <= 1'b1;
                  active_thread[(679*4)+2] <= 1'b1;
                  active_thread[(679*4)+3] <= 1'b1;
                  spc679_inst_done         <= `ARIANE_CORE679.piton_pc_vld;
                  spc679_phy_pc_w          <= `ARIANE_CORE679.piton_pc;
                end
            end
    

            assign spc680_thread_id = 2'b00;
            assign spc680_rtl_pc = spc680_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(680*4)]   <= 1'b0;
                  active_thread[(680*4)+1] <= 1'b0;
                  active_thread[(680*4)+2] <= 1'b0;
                  active_thread[(680*4)+3] <= 1'b0;
                  spc680_inst_done         <= 0;
                  spc680_phy_pc_w          <= 0;
                end else begin
                  active_thread[(680*4)]   <= 1'b1;
                  active_thread[(680*4)+1] <= 1'b1;
                  active_thread[(680*4)+2] <= 1'b1;
                  active_thread[(680*4)+3] <= 1'b1;
                  spc680_inst_done         <= `ARIANE_CORE680.piton_pc_vld;
                  spc680_phy_pc_w          <= `ARIANE_CORE680.piton_pc;
                end
            end
    

            assign spc681_thread_id = 2'b00;
            assign spc681_rtl_pc = spc681_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(681*4)]   <= 1'b0;
                  active_thread[(681*4)+1] <= 1'b0;
                  active_thread[(681*4)+2] <= 1'b0;
                  active_thread[(681*4)+3] <= 1'b0;
                  spc681_inst_done         <= 0;
                  spc681_phy_pc_w          <= 0;
                end else begin
                  active_thread[(681*4)]   <= 1'b1;
                  active_thread[(681*4)+1] <= 1'b1;
                  active_thread[(681*4)+2] <= 1'b1;
                  active_thread[(681*4)+3] <= 1'b1;
                  spc681_inst_done         <= `ARIANE_CORE681.piton_pc_vld;
                  spc681_phy_pc_w          <= `ARIANE_CORE681.piton_pc;
                end
            end
    

            assign spc682_thread_id = 2'b00;
            assign spc682_rtl_pc = spc682_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(682*4)]   <= 1'b0;
                  active_thread[(682*4)+1] <= 1'b0;
                  active_thread[(682*4)+2] <= 1'b0;
                  active_thread[(682*4)+3] <= 1'b0;
                  spc682_inst_done         <= 0;
                  spc682_phy_pc_w          <= 0;
                end else begin
                  active_thread[(682*4)]   <= 1'b1;
                  active_thread[(682*4)+1] <= 1'b1;
                  active_thread[(682*4)+2] <= 1'b1;
                  active_thread[(682*4)+3] <= 1'b1;
                  spc682_inst_done         <= `ARIANE_CORE682.piton_pc_vld;
                  spc682_phy_pc_w          <= `ARIANE_CORE682.piton_pc;
                end
            end
    

            assign spc683_thread_id = 2'b00;
            assign spc683_rtl_pc = spc683_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(683*4)]   <= 1'b0;
                  active_thread[(683*4)+1] <= 1'b0;
                  active_thread[(683*4)+2] <= 1'b0;
                  active_thread[(683*4)+3] <= 1'b0;
                  spc683_inst_done         <= 0;
                  spc683_phy_pc_w          <= 0;
                end else begin
                  active_thread[(683*4)]   <= 1'b1;
                  active_thread[(683*4)+1] <= 1'b1;
                  active_thread[(683*4)+2] <= 1'b1;
                  active_thread[(683*4)+3] <= 1'b1;
                  spc683_inst_done         <= `ARIANE_CORE683.piton_pc_vld;
                  spc683_phy_pc_w          <= `ARIANE_CORE683.piton_pc;
                end
            end
    

            assign spc684_thread_id = 2'b00;
            assign spc684_rtl_pc = spc684_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(684*4)]   <= 1'b0;
                  active_thread[(684*4)+1] <= 1'b0;
                  active_thread[(684*4)+2] <= 1'b0;
                  active_thread[(684*4)+3] <= 1'b0;
                  spc684_inst_done         <= 0;
                  spc684_phy_pc_w          <= 0;
                end else begin
                  active_thread[(684*4)]   <= 1'b1;
                  active_thread[(684*4)+1] <= 1'b1;
                  active_thread[(684*4)+2] <= 1'b1;
                  active_thread[(684*4)+3] <= 1'b1;
                  spc684_inst_done         <= `ARIANE_CORE684.piton_pc_vld;
                  spc684_phy_pc_w          <= `ARIANE_CORE684.piton_pc;
                end
            end
    

            assign spc685_thread_id = 2'b00;
            assign spc685_rtl_pc = spc685_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(685*4)]   <= 1'b0;
                  active_thread[(685*4)+1] <= 1'b0;
                  active_thread[(685*4)+2] <= 1'b0;
                  active_thread[(685*4)+3] <= 1'b0;
                  spc685_inst_done         <= 0;
                  spc685_phy_pc_w          <= 0;
                end else begin
                  active_thread[(685*4)]   <= 1'b1;
                  active_thread[(685*4)+1] <= 1'b1;
                  active_thread[(685*4)+2] <= 1'b1;
                  active_thread[(685*4)+3] <= 1'b1;
                  spc685_inst_done         <= `ARIANE_CORE685.piton_pc_vld;
                  spc685_phy_pc_w          <= `ARIANE_CORE685.piton_pc;
                end
            end
    

            assign spc686_thread_id = 2'b00;
            assign spc686_rtl_pc = spc686_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(686*4)]   <= 1'b0;
                  active_thread[(686*4)+1] <= 1'b0;
                  active_thread[(686*4)+2] <= 1'b0;
                  active_thread[(686*4)+3] <= 1'b0;
                  spc686_inst_done         <= 0;
                  spc686_phy_pc_w          <= 0;
                end else begin
                  active_thread[(686*4)]   <= 1'b1;
                  active_thread[(686*4)+1] <= 1'b1;
                  active_thread[(686*4)+2] <= 1'b1;
                  active_thread[(686*4)+3] <= 1'b1;
                  spc686_inst_done         <= `ARIANE_CORE686.piton_pc_vld;
                  spc686_phy_pc_w          <= `ARIANE_CORE686.piton_pc;
                end
            end
    

            assign spc687_thread_id = 2'b00;
            assign spc687_rtl_pc = spc687_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(687*4)]   <= 1'b0;
                  active_thread[(687*4)+1] <= 1'b0;
                  active_thread[(687*4)+2] <= 1'b0;
                  active_thread[(687*4)+3] <= 1'b0;
                  spc687_inst_done         <= 0;
                  spc687_phy_pc_w          <= 0;
                end else begin
                  active_thread[(687*4)]   <= 1'b1;
                  active_thread[(687*4)+1] <= 1'b1;
                  active_thread[(687*4)+2] <= 1'b1;
                  active_thread[(687*4)+3] <= 1'b1;
                  spc687_inst_done         <= `ARIANE_CORE687.piton_pc_vld;
                  spc687_phy_pc_w          <= `ARIANE_CORE687.piton_pc;
                end
            end
    

            assign spc688_thread_id = 2'b00;
            assign spc688_rtl_pc = spc688_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(688*4)]   <= 1'b0;
                  active_thread[(688*4)+1] <= 1'b0;
                  active_thread[(688*4)+2] <= 1'b0;
                  active_thread[(688*4)+3] <= 1'b0;
                  spc688_inst_done         <= 0;
                  spc688_phy_pc_w          <= 0;
                end else begin
                  active_thread[(688*4)]   <= 1'b1;
                  active_thread[(688*4)+1] <= 1'b1;
                  active_thread[(688*4)+2] <= 1'b1;
                  active_thread[(688*4)+3] <= 1'b1;
                  spc688_inst_done         <= `ARIANE_CORE688.piton_pc_vld;
                  spc688_phy_pc_w          <= `ARIANE_CORE688.piton_pc;
                end
            end
    

            assign spc689_thread_id = 2'b00;
            assign spc689_rtl_pc = spc689_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(689*4)]   <= 1'b0;
                  active_thread[(689*4)+1] <= 1'b0;
                  active_thread[(689*4)+2] <= 1'b0;
                  active_thread[(689*4)+3] <= 1'b0;
                  spc689_inst_done         <= 0;
                  spc689_phy_pc_w          <= 0;
                end else begin
                  active_thread[(689*4)]   <= 1'b1;
                  active_thread[(689*4)+1] <= 1'b1;
                  active_thread[(689*4)+2] <= 1'b1;
                  active_thread[(689*4)+3] <= 1'b1;
                  spc689_inst_done         <= `ARIANE_CORE689.piton_pc_vld;
                  spc689_phy_pc_w          <= `ARIANE_CORE689.piton_pc;
                end
            end
    

            assign spc690_thread_id = 2'b00;
            assign spc690_rtl_pc = spc690_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(690*4)]   <= 1'b0;
                  active_thread[(690*4)+1] <= 1'b0;
                  active_thread[(690*4)+2] <= 1'b0;
                  active_thread[(690*4)+3] <= 1'b0;
                  spc690_inst_done         <= 0;
                  spc690_phy_pc_w          <= 0;
                end else begin
                  active_thread[(690*4)]   <= 1'b1;
                  active_thread[(690*4)+1] <= 1'b1;
                  active_thread[(690*4)+2] <= 1'b1;
                  active_thread[(690*4)+3] <= 1'b1;
                  spc690_inst_done         <= `ARIANE_CORE690.piton_pc_vld;
                  spc690_phy_pc_w          <= `ARIANE_CORE690.piton_pc;
                end
            end
    

            assign spc691_thread_id = 2'b00;
            assign spc691_rtl_pc = spc691_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(691*4)]   <= 1'b0;
                  active_thread[(691*4)+1] <= 1'b0;
                  active_thread[(691*4)+2] <= 1'b0;
                  active_thread[(691*4)+3] <= 1'b0;
                  spc691_inst_done         <= 0;
                  spc691_phy_pc_w          <= 0;
                end else begin
                  active_thread[(691*4)]   <= 1'b1;
                  active_thread[(691*4)+1] <= 1'b1;
                  active_thread[(691*4)+2] <= 1'b1;
                  active_thread[(691*4)+3] <= 1'b1;
                  spc691_inst_done         <= `ARIANE_CORE691.piton_pc_vld;
                  spc691_phy_pc_w          <= `ARIANE_CORE691.piton_pc;
                end
            end
    

            assign spc692_thread_id = 2'b00;
            assign spc692_rtl_pc = spc692_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(692*4)]   <= 1'b0;
                  active_thread[(692*4)+1] <= 1'b0;
                  active_thread[(692*4)+2] <= 1'b0;
                  active_thread[(692*4)+3] <= 1'b0;
                  spc692_inst_done         <= 0;
                  spc692_phy_pc_w          <= 0;
                end else begin
                  active_thread[(692*4)]   <= 1'b1;
                  active_thread[(692*4)+1] <= 1'b1;
                  active_thread[(692*4)+2] <= 1'b1;
                  active_thread[(692*4)+3] <= 1'b1;
                  spc692_inst_done         <= `ARIANE_CORE692.piton_pc_vld;
                  spc692_phy_pc_w          <= `ARIANE_CORE692.piton_pc;
                end
            end
    

            assign spc693_thread_id = 2'b00;
            assign spc693_rtl_pc = spc693_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(693*4)]   <= 1'b0;
                  active_thread[(693*4)+1] <= 1'b0;
                  active_thread[(693*4)+2] <= 1'b0;
                  active_thread[(693*4)+3] <= 1'b0;
                  spc693_inst_done         <= 0;
                  spc693_phy_pc_w          <= 0;
                end else begin
                  active_thread[(693*4)]   <= 1'b1;
                  active_thread[(693*4)+1] <= 1'b1;
                  active_thread[(693*4)+2] <= 1'b1;
                  active_thread[(693*4)+3] <= 1'b1;
                  spc693_inst_done         <= `ARIANE_CORE693.piton_pc_vld;
                  spc693_phy_pc_w          <= `ARIANE_CORE693.piton_pc;
                end
            end
    

            assign spc694_thread_id = 2'b00;
            assign spc694_rtl_pc = spc694_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(694*4)]   <= 1'b0;
                  active_thread[(694*4)+1] <= 1'b0;
                  active_thread[(694*4)+2] <= 1'b0;
                  active_thread[(694*4)+3] <= 1'b0;
                  spc694_inst_done         <= 0;
                  spc694_phy_pc_w          <= 0;
                end else begin
                  active_thread[(694*4)]   <= 1'b1;
                  active_thread[(694*4)+1] <= 1'b1;
                  active_thread[(694*4)+2] <= 1'b1;
                  active_thread[(694*4)+3] <= 1'b1;
                  spc694_inst_done         <= `ARIANE_CORE694.piton_pc_vld;
                  spc694_phy_pc_w          <= `ARIANE_CORE694.piton_pc;
                end
            end
    

            assign spc695_thread_id = 2'b00;
            assign spc695_rtl_pc = spc695_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(695*4)]   <= 1'b0;
                  active_thread[(695*4)+1] <= 1'b0;
                  active_thread[(695*4)+2] <= 1'b0;
                  active_thread[(695*4)+3] <= 1'b0;
                  spc695_inst_done         <= 0;
                  spc695_phy_pc_w          <= 0;
                end else begin
                  active_thread[(695*4)]   <= 1'b1;
                  active_thread[(695*4)+1] <= 1'b1;
                  active_thread[(695*4)+2] <= 1'b1;
                  active_thread[(695*4)+3] <= 1'b1;
                  spc695_inst_done         <= `ARIANE_CORE695.piton_pc_vld;
                  spc695_phy_pc_w          <= `ARIANE_CORE695.piton_pc;
                end
            end
    

            assign spc696_thread_id = 2'b00;
            assign spc696_rtl_pc = spc696_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(696*4)]   <= 1'b0;
                  active_thread[(696*4)+1] <= 1'b0;
                  active_thread[(696*4)+2] <= 1'b0;
                  active_thread[(696*4)+3] <= 1'b0;
                  spc696_inst_done         <= 0;
                  spc696_phy_pc_w          <= 0;
                end else begin
                  active_thread[(696*4)]   <= 1'b1;
                  active_thread[(696*4)+1] <= 1'b1;
                  active_thread[(696*4)+2] <= 1'b1;
                  active_thread[(696*4)+3] <= 1'b1;
                  spc696_inst_done         <= `ARIANE_CORE696.piton_pc_vld;
                  spc696_phy_pc_w          <= `ARIANE_CORE696.piton_pc;
                end
            end
    

            assign spc697_thread_id = 2'b00;
            assign spc697_rtl_pc = spc697_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(697*4)]   <= 1'b0;
                  active_thread[(697*4)+1] <= 1'b0;
                  active_thread[(697*4)+2] <= 1'b0;
                  active_thread[(697*4)+3] <= 1'b0;
                  spc697_inst_done         <= 0;
                  spc697_phy_pc_w          <= 0;
                end else begin
                  active_thread[(697*4)]   <= 1'b1;
                  active_thread[(697*4)+1] <= 1'b1;
                  active_thread[(697*4)+2] <= 1'b1;
                  active_thread[(697*4)+3] <= 1'b1;
                  spc697_inst_done         <= `ARIANE_CORE697.piton_pc_vld;
                  spc697_phy_pc_w          <= `ARIANE_CORE697.piton_pc;
                end
            end
    

            assign spc698_thread_id = 2'b00;
            assign spc698_rtl_pc = spc698_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(698*4)]   <= 1'b0;
                  active_thread[(698*4)+1] <= 1'b0;
                  active_thread[(698*4)+2] <= 1'b0;
                  active_thread[(698*4)+3] <= 1'b0;
                  spc698_inst_done         <= 0;
                  spc698_phy_pc_w          <= 0;
                end else begin
                  active_thread[(698*4)]   <= 1'b1;
                  active_thread[(698*4)+1] <= 1'b1;
                  active_thread[(698*4)+2] <= 1'b1;
                  active_thread[(698*4)+3] <= 1'b1;
                  spc698_inst_done         <= `ARIANE_CORE698.piton_pc_vld;
                  spc698_phy_pc_w          <= `ARIANE_CORE698.piton_pc;
                end
            end
    

            assign spc699_thread_id = 2'b00;
            assign spc699_rtl_pc = spc699_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(699*4)]   <= 1'b0;
                  active_thread[(699*4)+1] <= 1'b0;
                  active_thread[(699*4)+2] <= 1'b0;
                  active_thread[(699*4)+3] <= 1'b0;
                  spc699_inst_done         <= 0;
                  spc699_phy_pc_w          <= 0;
                end else begin
                  active_thread[(699*4)]   <= 1'b1;
                  active_thread[(699*4)+1] <= 1'b1;
                  active_thread[(699*4)+2] <= 1'b1;
                  active_thread[(699*4)+3] <= 1'b1;
                  spc699_inst_done         <= `ARIANE_CORE699.piton_pc_vld;
                  spc699_phy_pc_w          <= `ARIANE_CORE699.piton_pc;
                end
            end
    

            assign spc700_thread_id = 2'b00;
            assign spc700_rtl_pc = spc700_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(700*4)]   <= 1'b0;
                  active_thread[(700*4)+1] <= 1'b0;
                  active_thread[(700*4)+2] <= 1'b0;
                  active_thread[(700*4)+3] <= 1'b0;
                  spc700_inst_done         <= 0;
                  spc700_phy_pc_w          <= 0;
                end else begin
                  active_thread[(700*4)]   <= 1'b1;
                  active_thread[(700*4)+1] <= 1'b1;
                  active_thread[(700*4)+2] <= 1'b1;
                  active_thread[(700*4)+3] <= 1'b1;
                  spc700_inst_done         <= `ARIANE_CORE700.piton_pc_vld;
                  spc700_phy_pc_w          <= `ARIANE_CORE700.piton_pc;
                end
            end
    

            assign spc701_thread_id = 2'b00;
            assign spc701_rtl_pc = spc701_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(701*4)]   <= 1'b0;
                  active_thread[(701*4)+1] <= 1'b0;
                  active_thread[(701*4)+2] <= 1'b0;
                  active_thread[(701*4)+3] <= 1'b0;
                  spc701_inst_done         <= 0;
                  spc701_phy_pc_w          <= 0;
                end else begin
                  active_thread[(701*4)]   <= 1'b1;
                  active_thread[(701*4)+1] <= 1'b1;
                  active_thread[(701*4)+2] <= 1'b1;
                  active_thread[(701*4)+3] <= 1'b1;
                  spc701_inst_done         <= `ARIANE_CORE701.piton_pc_vld;
                  spc701_phy_pc_w          <= `ARIANE_CORE701.piton_pc;
                end
            end
    

            assign spc702_thread_id = 2'b00;
            assign spc702_rtl_pc = spc702_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(702*4)]   <= 1'b0;
                  active_thread[(702*4)+1] <= 1'b0;
                  active_thread[(702*4)+2] <= 1'b0;
                  active_thread[(702*4)+3] <= 1'b0;
                  spc702_inst_done         <= 0;
                  spc702_phy_pc_w          <= 0;
                end else begin
                  active_thread[(702*4)]   <= 1'b1;
                  active_thread[(702*4)+1] <= 1'b1;
                  active_thread[(702*4)+2] <= 1'b1;
                  active_thread[(702*4)+3] <= 1'b1;
                  spc702_inst_done         <= `ARIANE_CORE702.piton_pc_vld;
                  spc702_phy_pc_w          <= `ARIANE_CORE702.piton_pc;
                end
            end
    

            assign spc703_thread_id = 2'b00;
            assign spc703_rtl_pc = spc703_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(703*4)]   <= 1'b0;
                  active_thread[(703*4)+1] <= 1'b0;
                  active_thread[(703*4)+2] <= 1'b0;
                  active_thread[(703*4)+3] <= 1'b0;
                  spc703_inst_done         <= 0;
                  spc703_phy_pc_w          <= 0;
                end else begin
                  active_thread[(703*4)]   <= 1'b1;
                  active_thread[(703*4)+1] <= 1'b1;
                  active_thread[(703*4)+2] <= 1'b1;
                  active_thread[(703*4)+3] <= 1'b1;
                  spc703_inst_done         <= `ARIANE_CORE703.piton_pc_vld;
                  spc703_phy_pc_w          <= `ARIANE_CORE703.piton_pc;
                end
            end
    

            assign spc704_thread_id = 2'b00;
            assign spc704_rtl_pc = spc704_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(704*4)]   <= 1'b0;
                  active_thread[(704*4)+1] <= 1'b0;
                  active_thread[(704*4)+2] <= 1'b0;
                  active_thread[(704*4)+3] <= 1'b0;
                  spc704_inst_done         <= 0;
                  spc704_phy_pc_w          <= 0;
                end else begin
                  active_thread[(704*4)]   <= 1'b1;
                  active_thread[(704*4)+1] <= 1'b1;
                  active_thread[(704*4)+2] <= 1'b1;
                  active_thread[(704*4)+3] <= 1'b1;
                  spc704_inst_done         <= `ARIANE_CORE704.piton_pc_vld;
                  spc704_phy_pc_w          <= `ARIANE_CORE704.piton_pc;
                end
            end
    

            assign spc705_thread_id = 2'b00;
            assign spc705_rtl_pc = spc705_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(705*4)]   <= 1'b0;
                  active_thread[(705*4)+1] <= 1'b0;
                  active_thread[(705*4)+2] <= 1'b0;
                  active_thread[(705*4)+3] <= 1'b0;
                  spc705_inst_done         <= 0;
                  spc705_phy_pc_w          <= 0;
                end else begin
                  active_thread[(705*4)]   <= 1'b1;
                  active_thread[(705*4)+1] <= 1'b1;
                  active_thread[(705*4)+2] <= 1'b1;
                  active_thread[(705*4)+3] <= 1'b1;
                  spc705_inst_done         <= `ARIANE_CORE705.piton_pc_vld;
                  spc705_phy_pc_w          <= `ARIANE_CORE705.piton_pc;
                end
            end
    

            assign spc706_thread_id = 2'b00;
            assign spc706_rtl_pc = spc706_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(706*4)]   <= 1'b0;
                  active_thread[(706*4)+1] <= 1'b0;
                  active_thread[(706*4)+2] <= 1'b0;
                  active_thread[(706*4)+3] <= 1'b0;
                  spc706_inst_done         <= 0;
                  spc706_phy_pc_w          <= 0;
                end else begin
                  active_thread[(706*4)]   <= 1'b1;
                  active_thread[(706*4)+1] <= 1'b1;
                  active_thread[(706*4)+2] <= 1'b1;
                  active_thread[(706*4)+3] <= 1'b1;
                  spc706_inst_done         <= `ARIANE_CORE706.piton_pc_vld;
                  spc706_phy_pc_w          <= `ARIANE_CORE706.piton_pc;
                end
            end
    

            assign spc707_thread_id = 2'b00;
            assign spc707_rtl_pc = spc707_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(707*4)]   <= 1'b0;
                  active_thread[(707*4)+1] <= 1'b0;
                  active_thread[(707*4)+2] <= 1'b0;
                  active_thread[(707*4)+3] <= 1'b0;
                  spc707_inst_done         <= 0;
                  spc707_phy_pc_w          <= 0;
                end else begin
                  active_thread[(707*4)]   <= 1'b1;
                  active_thread[(707*4)+1] <= 1'b1;
                  active_thread[(707*4)+2] <= 1'b1;
                  active_thread[(707*4)+3] <= 1'b1;
                  spc707_inst_done         <= `ARIANE_CORE707.piton_pc_vld;
                  spc707_phy_pc_w          <= `ARIANE_CORE707.piton_pc;
                end
            end
    

            assign spc708_thread_id = 2'b00;
            assign spc708_rtl_pc = spc708_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(708*4)]   <= 1'b0;
                  active_thread[(708*4)+1] <= 1'b0;
                  active_thread[(708*4)+2] <= 1'b0;
                  active_thread[(708*4)+3] <= 1'b0;
                  spc708_inst_done         <= 0;
                  spc708_phy_pc_w          <= 0;
                end else begin
                  active_thread[(708*4)]   <= 1'b1;
                  active_thread[(708*4)+1] <= 1'b1;
                  active_thread[(708*4)+2] <= 1'b1;
                  active_thread[(708*4)+3] <= 1'b1;
                  spc708_inst_done         <= `ARIANE_CORE708.piton_pc_vld;
                  spc708_phy_pc_w          <= `ARIANE_CORE708.piton_pc;
                end
            end
    

            assign spc709_thread_id = 2'b00;
            assign spc709_rtl_pc = spc709_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(709*4)]   <= 1'b0;
                  active_thread[(709*4)+1] <= 1'b0;
                  active_thread[(709*4)+2] <= 1'b0;
                  active_thread[(709*4)+3] <= 1'b0;
                  spc709_inst_done         <= 0;
                  spc709_phy_pc_w          <= 0;
                end else begin
                  active_thread[(709*4)]   <= 1'b1;
                  active_thread[(709*4)+1] <= 1'b1;
                  active_thread[(709*4)+2] <= 1'b1;
                  active_thread[(709*4)+3] <= 1'b1;
                  spc709_inst_done         <= `ARIANE_CORE709.piton_pc_vld;
                  spc709_phy_pc_w          <= `ARIANE_CORE709.piton_pc;
                end
            end
    

            assign spc710_thread_id = 2'b00;
            assign spc710_rtl_pc = spc710_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(710*4)]   <= 1'b0;
                  active_thread[(710*4)+1] <= 1'b0;
                  active_thread[(710*4)+2] <= 1'b0;
                  active_thread[(710*4)+3] <= 1'b0;
                  spc710_inst_done         <= 0;
                  spc710_phy_pc_w          <= 0;
                end else begin
                  active_thread[(710*4)]   <= 1'b1;
                  active_thread[(710*4)+1] <= 1'b1;
                  active_thread[(710*4)+2] <= 1'b1;
                  active_thread[(710*4)+3] <= 1'b1;
                  spc710_inst_done         <= `ARIANE_CORE710.piton_pc_vld;
                  spc710_phy_pc_w          <= `ARIANE_CORE710.piton_pc;
                end
            end
    

            assign spc711_thread_id = 2'b00;
            assign spc711_rtl_pc = spc711_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(711*4)]   <= 1'b0;
                  active_thread[(711*4)+1] <= 1'b0;
                  active_thread[(711*4)+2] <= 1'b0;
                  active_thread[(711*4)+3] <= 1'b0;
                  spc711_inst_done         <= 0;
                  spc711_phy_pc_w          <= 0;
                end else begin
                  active_thread[(711*4)]   <= 1'b1;
                  active_thread[(711*4)+1] <= 1'b1;
                  active_thread[(711*4)+2] <= 1'b1;
                  active_thread[(711*4)+3] <= 1'b1;
                  spc711_inst_done         <= `ARIANE_CORE711.piton_pc_vld;
                  spc711_phy_pc_w          <= `ARIANE_CORE711.piton_pc;
                end
            end
    

            assign spc712_thread_id = 2'b00;
            assign spc712_rtl_pc = spc712_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(712*4)]   <= 1'b0;
                  active_thread[(712*4)+1] <= 1'b0;
                  active_thread[(712*4)+2] <= 1'b0;
                  active_thread[(712*4)+3] <= 1'b0;
                  spc712_inst_done         <= 0;
                  spc712_phy_pc_w          <= 0;
                end else begin
                  active_thread[(712*4)]   <= 1'b1;
                  active_thread[(712*4)+1] <= 1'b1;
                  active_thread[(712*4)+2] <= 1'b1;
                  active_thread[(712*4)+3] <= 1'b1;
                  spc712_inst_done         <= `ARIANE_CORE712.piton_pc_vld;
                  spc712_phy_pc_w          <= `ARIANE_CORE712.piton_pc;
                end
            end
    

            assign spc713_thread_id = 2'b00;
            assign spc713_rtl_pc = spc713_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(713*4)]   <= 1'b0;
                  active_thread[(713*4)+1] <= 1'b0;
                  active_thread[(713*4)+2] <= 1'b0;
                  active_thread[(713*4)+3] <= 1'b0;
                  spc713_inst_done         <= 0;
                  spc713_phy_pc_w          <= 0;
                end else begin
                  active_thread[(713*4)]   <= 1'b1;
                  active_thread[(713*4)+1] <= 1'b1;
                  active_thread[(713*4)+2] <= 1'b1;
                  active_thread[(713*4)+3] <= 1'b1;
                  spc713_inst_done         <= `ARIANE_CORE713.piton_pc_vld;
                  spc713_phy_pc_w          <= `ARIANE_CORE713.piton_pc;
                end
            end
    

            assign spc714_thread_id = 2'b00;
            assign spc714_rtl_pc = spc714_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(714*4)]   <= 1'b0;
                  active_thread[(714*4)+1] <= 1'b0;
                  active_thread[(714*4)+2] <= 1'b0;
                  active_thread[(714*4)+3] <= 1'b0;
                  spc714_inst_done         <= 0;
                  spc714_phy_pc_w          <= 0;
                end else begin
                  active_thread[(714*4)]   <= 1'b1;
                  active_thread[(714*4)+1] <= 1'b1;
                  active_thread[(714*4)+2] <= 1'b1;
                  active_thread[(714*4)+3] <= 1'b1;
                  spc714_inst_done         <= `ARIANE_CORE714.piton_pc_vld;
                  spc714_phy_pc_w          <= `ARIANE_CORE714.piton_pc;
                end
            end
    

            assign spc715_thread_id = 2'b00;
            assign spc715_rtl_pc = spc715_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(715*4)]   <= 1'b0;
                  active_thread[(715*4)+1] <= 1'b0;
                  active_thread[(715*4)+2] <= 1'b0;
                  active_thread[(715*4)+3] <= 1'b0;
                  spc715_inst_done         <= 0;
                  spc715_phy_pc_w          <= 0;
                end else begin
                  active_thread[(715*4)]   <= 1'b1;
                  active_thread[(715*4)+1] <= 1'b1;
                  active_thread[(715*4)+2] <= 1'b1;
                  active_thread[(715*4)+3] <= 1'b1;
                  spc715_inst_done         <= `ARIANE_CORE715.piton_pc_vld;
                  spc715_phy_pc_w          <= `ARIANE_CORE715.piton_pc;
                end
            end
    

            assign spc716_thread_id = 2'b00;
            assign spc716_rtl_pc = spc716_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(716*4)]   <= 1'b0;
                  active_thread[(716*4)+1] <= 1'b0;
                  active_thread[(716*4)+2] <= 1'b0;
                  active_thread[(716*4)+3] <= 1'b0;
                  spc716_inst_done         <= 0;
                  spc716_phy_pc_w          <= 0;
                end else begin
                  active_thread[(716*4)]   <= 1'b1;
                  active_thread[(716*4)+1] <= 1'b1;
                  active_thread[(716*4)+2] <= 1'b1;
                  active_thread[(716*4)+3] <= 1'b1;
                  spc716_inst_done         <= `ARIANE_CORE716.piton_pc_vld;
                  spc716_phy_pc_w          <= `ARIANE_CORE716.piton_pc;
                end
            end
    

            assign spc717_thread_id = 2'b00;
            assign spc717_rtl_pc = spc717_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(717*4)]   <= 1'b0;
                  active_thread[(717*4)+1] <= 1'b0;
                  active_thread[(717*4)+2] <= 1'b0;
                  active_thread[(717*4)+3] <= 1'b0;
                  spc717_inst_done         <= 0;
                  spc717_phy_pc_w          <= 0;
                end else begin
                  active_thread[(717*4)]   <= 1'b1;
                  active_thread[(717*4)+1] <= 1'b1;
                  active_thread[(717*4)+2] <= 1'b1;
                  active_thread[(717*4)+3] <= 1'b1;
                  spc717_inst_done         <= `ARIANE_CORE717.piton_pc_vld;
                  spc717_phy_pc_w          <= `ARIANE_CORE717.piton_pc;
                end
            end
    

            assign spc718_thread_id = 2'b00;
            assign spc718_rtl_pc = spc718_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(718*4)]   <= 1'b0;
                  active_thread[(718*4)+1] <= 1'b0;
                  active_thread[(718*4)+2] <= 1'b0;
                  active_thread[(718*4)+3] <= 1'b0;
                  spc718_inst_done         <= 0;
                  spc718_phy_pc_w          <= 0;
                end else begin
                  active_thread[(718*4)]   <= 1'b1;
                  active_thread[(718*4)+1] <= 1'b1;
                  active_thread[(718*4)+2] <= 1'b1;
                  active_thread[(718*4)+3] <= 1'b1;
                  spc718_inst_done         <= `ARIANE_CORE718.piton_pc_vld;
                  spc718_phy_pc_w          <= `ARIANE_CORE718.piton_pc;
                end
            end
    

            assign spc719_thread_id = 2'b00;
            assign spc719_rtl_pc = spc719_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(719*4)]   <= 1'b0;
                  active_thread[(719*4)+1] <= 1'b0;
                  active_thread[(719*4)+2] <= 1'b0;
                  active_thread[(719*4)+3] <= 1'b0;
                  spc719_inst_done         <= 0;
                  spc719_phy_pc_w          <= 0;
                end else begin
                  active_thread[(719*4)]   <= 1'b1;
                  active_thread[(719*4)+1] <= 1'b1;
                  active_thread[(719*4)+2] <= 1'b1;
                  active_thread[(719*4)+3] <= 1'b1;
                  spc719_inst_done         <= `ARIANE_CORE719.piton_pc_vld;
                  spc719_phy_pc_w          <= `ARIANE_CORE719.piton_pc;
                end
            end
    

            assign spc720_thread_id = 2'b00;
            assign spc720_rtl_pc = spc720_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(720*4)]   <= 1'b0;
                  active_thread[(720*4)+1] <= 1'b0;
                  active_thread[(720*4)+2] <= 1'b0;
                  active_thread[(720*4)+3] <= 1'b0;
                  spc720_inst_done         <= 0;
                  spc720_phy_pc_w          <= 0;
                end else begin
                  active_thread[(720*4)]   <= 1'b1;
                  active_thread[(720*4)+1] <= 1'b1;
                  active_thread[(720*4)+2] <= 1'b1;
                  active_thread[(720*4)+3] <= 1'b1;
                  spc720_inst_done         <= `ARIANE_CORE720.piton_pc_vld;
                  spc720_phy_pc_w          <= `ARIANE_CORE720.piton_pc;
                end
            end
    

            assign spc721_thread_id = 2'b00;
            assign spc721_rtl_pc = spc721_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(721*4)]   <= 1'b0;
                  active_thread[(721*4)+1] <= 1'b0;
                  active_thread[(721*4)+2] <= 1'b0;
                  active_thread[(721*4)+3] <= 1'b0;
                  spc721_inst_done         <= 0;
                  spc721_phy_pc_w          <= 0;
                end else begin
                  active_thread[(721*4)]   <= 1'b1;
                  active_thread[(721*4)+1] <= 1'b1;
                  active_thread[(721*4)+2] <= 1'b1;
                  active_thread[(721*4)+3] <= 1'b1;
                  spc721_inst_done         <= `ARIANE_CORE721.piton_pc_vld;
                  spc721_phy_pc_w          <= `ARIANE_CORE721.piton_pc;
                end
            end
    

            assign spc722_thread_id = 2'b00;
            assign spc722_rtl_pc = spc722_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(722*4)]   <= 1'b0;
                  active_thread[(722*4)+1] <= 1'b0;
                  active_thread[(722*4)+2] <= 1'b0;
                  active_thread[(722*4)+3] <= 1'b0;
                  spc722_inst_done         <= 0;
                  spc722_phy_pc_w          <= 0;
                end else begin
                  active_thread[(722*4)]   <= 1'b1;
                  active_thread[(722*4)+1] <= 1'b1;
                  active_thread[(722*4)+2] <= 1'b1;
                  active_thread[(722*4)+3] <= 1'b1;
                  spc722_inst_done         <= `ARIANE_CORE722.piton_pc_vld;
                  spc722_phy_pc_w          <= `ARIANE_CORE722.piton_pc;
                end
            end
    

            assign spc723_thread_id = 2'b00;
            assign spc723_rtl_pc = spc723_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(723*4)]   <= 1'b0;
                  active_thread[(723*4)+1] <= 1'b0;
                  active_thread[(723*4)+2] <= 1'b0;
                  active_thread[(723*4)+3] <= 1'b0;
                  spc723_inst_done         <= 0;
                  spc723_phy_pc_w          <= 0;
                end else begin
                  active_thread[(723*4)]   <= 1'b1;
                  active_thread[(723*4)+1] <= 1'b1;
                  active_thread[(723*4)+2] <= 1'b1;
                  active_thread[(723*4)+3] <= 1'b1;
                  spc723_inst_done         <= `ARIANE_CORE723.piton_pc_vld;
                  spc723_phy_pc_w          <= `ARIANE_CORE723.piton_pc;
                end
            end
    

            assign spc724_thread_id = 2'b00;
            assign spc724_rtl_pc = spc724_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(724*4)]   <= 1'b0;
                  active_thread[(724*4)+1] <= 1'b0;
                  active_thread[(724*4)+2] <= 1'b0;
                  active_thread[(724*4)+3] <= 1'b0;
                  spc724_inst_done         <= 0;
                  spc724_phy_pc_w          <= 0;
                end else begin
                  active_thread[(724*4)]   <= 1'b1;
                  active_thread[(724*4)+1] <= 1'b1;
                  active_thread[(724*4)+2] <= 1'b1;
                  active_thread[(724*4)+3] <= 1'b1;
                  spc724_inst_done         <= `ARIANE_CORE724.piton_pc_vld;
                  spc724_phy_pc_w          <= `ARIANE_CORE724.piton_pc;
                end
            end
    

            assign spc725_thread_id = 2'b00;
            assign spc725_rtl_pc = spc725_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(725*4)]   <= 1'b0;
                  active_thread[(725*4)+1] <= 1'b0;
                  active_thread[(725*4)+2] <= 1'b0;
                  active_thread[(725*4)+3] <= 1'b0;
                  spc725_inst_done         <= 0;
                  spc725_phy_pc_w          <= 0;
                end else begin
                  active_thread[(725*4)]   <= 1'b1;
                  active_thread[(725*4)+1] <= 1'b1;
                  active_thread[(725*4)+2] <= 1'b1;
                  active_thread[(725*4)+3] <= 1'b1;
                  spc725_inst_done         <= `ARIANE_CORE725.piton_pc_vld;
                  spc725_phy_pc_w          <= `ARIANE_CORE725.piton_pc;
                end
            end
    

            assign spc726_thread_id = 2'b00;
            assign spc726_rtl_pc = spc726_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(726*4)]   <= 1'b0;
                  active_thread[(726*4)+1] <= 1'b0;
                  active_thread[(726*4)+2] <= 1'b0;
                  active_thread[(726*4)+3] <= 1'b0;
                  spc726_inst_done         <= 0;
                  spc726_phy_pc_w          <= 0;
                end else begin
                  active_thread[(726*4)]   <= 1'b1;
                  active_thread[(726*4)+1] <= 1'b1;
                  active_thread[(726*4)+2] <= 1'b1;
                  active_thread[(726*4)+3] <= 1'b1;
                  spc726_inst_done         <= `ARIANE_CORE726.piton_pc_vld;
                  spc726_phy_pc_w          <= `ARIANE_CORE726.piton_pc;
                end
            end
    

            assign spc727_thread_id = 2'b00;
            assign spc727_rtl_pc = spc727_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(727*4)]   <= 1'b0;
                  active_thread[(727*4)+1] <= 1'b0;
                  active_thread[(727*4)+2] <= 1'b0;
                  active_thread[(727*4)+3] <= 1'b0;
                  spc727_inst_done         <= 0;
                  spc727_phy_pc_w          <= 0;
                end else begin
                  active_thread[(727*4)]   <= 1'b1;
                  active_thread[(727*4)+1] <= 1'b1;
                  active_thread[(727*4)+2] <= 1'b1;
                  active_thread[(727*4)+3] <= 1'b1;
                  spc727_inst_done         <= `ARIANE_CORE727.piton_pc_vld;
                  spc727_phy_pc_w          <= `ARIANE_CORE727.piton_pc;
                end
            end
    

            assign spc728_thread_id = 2'b00;
            assign spc728_rtl_pc = spc728_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(728*4)]   <= 1'b0;
                  active_thread[(728*4)+1] <= 1'b0;
                  active_thread[(728*4)+2] <= 1'b0;
                  active_thread[(728*4)+3] <= 1'b0;
                  spc728_inst_done         <= 0;
                  spc728_phy_pc_w          <= 0;
                end else begin
                  active_thread[(728*4)]   <= 1'b1;
                  active_thread[(728*4)+1] <= 1'b1;
                  active_thread[(728*4)+2] <= 1'b1;
                  active_thread[(728*4)+3] <= 1'b1;
                  spc728_inst_done         <= `ARIANE_CORE728.piton_pc_vld;
                  spc728_phy_pc_w          <= `ARIANE_CORE728.piton_pc;
                end
            end
    

            assign spc729_thread_id = 2'b00;
            assign spc729_rtl_pc = spc729_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(729*4)]   <= 1'b0;
                  active_thread[(729*4)+1] <= 1'b0;
                  active_thread[(729*4)+2] <= 1'b0;
                  active_thread[(729*4)+3] <= 1'b0;
                  spc729_inst_done         <= 0;
                  spc729_phy_pc_w          <= 0;
                end else begin
                  active_thread[(729*4)]   <= 1'b1;
                  active_thread[(729*4)+1] <= 1'b1;
                  active_thread[(729*4)+2] <= 1'b1;
                  active_thread[(729*4)+3] <= 1'b1;
                  spc729_inst_done         <= `ARIANE_CORE729.piton_pc_vld;
                  spc729_phy_pc_w          <= `ARIANE_CORE729.piton_pc;
                end
            end
    

            assign spc730_thread_id = 2'b00;
            assign spc730_rtl_pc = spc730_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(730*4)]   <= 1'b0;
                  active_thread[(730*4)+1] <= 1'b0;
                  active_thread[(730*4)+2] <= 1'b0;
                  active_thread[(730*4)+3] <= 1'b0;
                  spc730_inst_done         <= 0;
                  spc730_phy_pc_w          <= 0;
                end else begin
                  active_thread[(730*4)]   <= 1'b1;
                  active_thread[(730*4)+1] <= 1'b1;
                  active_thread[(730*4)+2] <= 1'b1;
                  active_thread[(730*4)+3] <= 1'b1;
                  spc730_inst_done         <= `ARIANE_CORE730.piton_pc_vld;
                  spc730_phy_pc_w          <= `ARIANE_CORE730.piton_pc;
                end
            end
    

            assign spc731_thread_id = 2'b00;
            assign spc731_rtl_pc = spc731_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(731*4)]   <= 1'b0;
                  active_thread[(731*4)+1] <= 1'b0;
                  active_thread[(731*4)+2] <= 1'b0;
                  active_thread[(731*4)+3] <= 1'b0;
                  spc731_inst_done         <= 0;
                  spc731_phy_pc_w          <= 0;
                end else begin
                  active_thread[(731*4)]   <= 1'b1;
                  active_thread[(731*4)+1] <= 1'b1;
                  active_thread[(731*4)+2] <= 1'b1;
                  active_thread[(731*4)+3] <= 1'b1;
                  spc731_inst_done         <= `ARIANE_CORE731.piton_pc_vld;
                  spc731_phy_pc_w          <= `ARIANE_CORE731.piton_pc;
                end
            end
    

            assign spc732_thread_id = 2'b00;
            assign spc732_rtl_pc = spc732_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(732*4)]   <= 1'b0;
                  active_thread[(732*4)+1] <= 1'b0;
                  active_thread[(732*4)+2] <= 1'b0;
                  active_thread[(732*4)+3] <= 1'b0;
                  spc732_inst_done         <= 0;
                  spc732_phy_pc_w          <= 0;
                end else begin
                  active_thread[(732*4)]   <= 1'b1;
                  active_thread[(732*4)+1] <= 1'b1;
                  active_thread[(732*4)+2] <= 1'b1;
                  active_thread[(732*4)+3] <= 1'b1;
                  spc732_inst_done         <= `ARIANE_CORE732.piton_pc_vld;
                  spc732_phy_pc_w          <= `ARIANE_CORE732.piton_pc;
                end
            end
    

            assign spc733_thread_id = 2'b00;
            assign spc733_rtl_pc = spc733_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(733*4)]   <= 1'b0;
                  active_thread[(733*4)+1] <= 1'b0;
                  active_thread[(733*4)+2] <= 1'b0;
                  active_thread[(733*4)+3] <= 1'b0;
                  spc733_inst_done         <= 0;
                  spc733_phy_pc_w          <= 0;
                end else begin
                  active_thread[(733*4)]   <= 1'b1;
                  active_thread[(733*4)+1] <= 1'b1;
                  active_thread[(733*4)+2] <= 1'b1;
                  active_thread[(733*4)+3] <= 1'b1;
                  spc733_inst_done         <= `ARIANE_CORE733.piton_pc_vld;
                  spc733_phy_pc_w          <= `ARIANE_CORE733.piton_pc;
                end
            end
    

            assign spc734_thread_id = 2'b00;
            assign spc734_rtl_pc = spc734_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(734*4)]   <= 1'b0;
                  active_thread[(734*4)+1] <= 1'b0;
                  active_thread[(734*4)+2] <= 1'b0;
                  active_thread[(734*4)+3] <= 1'b0;
                  spc734_inst_done         <= 0;
                  spc734_phy_pc_w          <= 0;
                end else begin
                  active_thread[(734*4)]   <= 1'b1;
                  active_thread[(734*4)+1] <= 1'b1;
                  active_thread[(734*4)+2] <= 1'b1;
                  active_thread[(734*4)+3] <= 1'b1;
                  spc734_inst_done         <= `ARIANE_CORE734.piton_pc_vld;
                  spc734_phy_pc_w          <= `ARIANE_CORE734.piton_pc;
                end
            end
    

            assign spc735_thread_id = 2'b00;
            assign spc735_rtl_pc = spc735_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(735*4)]   <= 1'b0;
                  active_thread[(735*4)+1] <= 1'b0;
                  active_thread[(735*4)+2] <= 1'b0;
                  active_thread[(735*4)+3] <= 1'b0;
                  spc735_inst_done         <= 0;
                  spc735_phy_pc_w          <= 0;
                end else begin
                  active_thread[(735*4)]   <= 1'b1;
                  active_thread[(735*4)+1] <= 1'b1;
                  active_thread[(735*4)+2] <= 1'b1;
                  active_thread[(735*4)+3] <= 1'b1;
                  spc735_inst_done         <= `ARIANE_CORE735.piton_pc_vld;
                  spc735_phy_pc_w          <= `ARIANE_CORE735.piton_pc;
                end
            end
    

            assign spc736_thread_id = 2'b00;
            assign spc736_rtl_pc = spc736_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(736*4)]   <= 1'b0;
                  active_thread[(736*4)+1] <= 1'b0;
                  active_thread[(736*4)+2] <= 1'b0;
                  active_thread[(736*4)+3] <= 1'b0;
                  spc736_inst_done         <= 0;
                  spc736_phy_pc_w          <= 0;
                end else begin
                  active_thread[(736*4)]   <= 1'b1;
                  active_thread[(736*4)+1] <= 1'b1;
                  active_thread[(736*4)+2] <= 1'b1;
                  active_thread[(736*4)+3] <= 1'b1;
                  spc736_inst_done         <= `ARIANE_CORE736.piton_pc_vld;
                  spc736_phy_pc_w          <= `ARIANE_CORE736.piton_pc;
                end
            end
    

            assign spc737_thread_id = 2'b00;
            assign spc737_rtl_pc = spc737_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(737*4)]   <= 1'b0;
                  active_thread[(737*4)+1] <= 1'b0;
                  active_thread[(737*4)+2] <= 1'b0;
                  active_thread[(737*4)+3] <= 1'b0;
                  spc737_inst_done         <= 0;
                  spc737_phy_pc_w          <= 0;
                end else begin
                  active_thread[(737*4)]   <= 1'b1;
                  active_thread[(737*4)+1] <= 1'b1;
                  active_thread[(737*4)+2] <= 1'b1;
                  active_thread[(737*4)+3] <= 1'b1;
                  spc737_inst_done         <= `ARIANE_CORE737.piton_pc_vld;
                  spc737_phy_pc_w          <= `ARIANE_CORE737.piton_pc;
                end
            end
    

            assign spc738_thread_id = 2'b00;
            assign spc738_rtl_pc = spc738_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(738*4)]   <= 1'b0;
                  active_thread[(738*4)+1] <= 1'b0;
                  active_thread[(738*4)+2] <= 1'b0;
                  active_thread[(738*4)+3] <= 1'b0;
                  spc738_inst_done         <= 0;
                  spc738_phy_pc_w          <= 0;
                end else begin
                  active_thread[(738*4)]   <= 1'b1;
                  active_thread[(738*4)+1] <= 1'b1;
                  active_thread[(738*4)+2] <= 1'b1;
                  active_thread[(738*4)+3] <= 1'b1;
                  spc738_inst_done         <= `ARIANE_CORE738.piton_pc_vld;
                  spc738_phy_pc_w          <= `ARIANE_CORE738.piton_pc;
                end
            end
    

            assign spc739_thread_id = 2'b00;
            assign spc739_rtl_pc = spc739_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(739*4)]   <= 1'b0;
                  active_thread[(739*4)+1] <= 1'b0;
                  active_thread[(739*4)+2] <= 1'b0;
                  active_thread[(739*4)+3] <= 1'b0;
                  spc739_inst_done         <= 0;
                  spc739_phy_pc_w          <= 0;
                end else begin
                  active_thread[(739*4)]   <= 1'b1;
                  active_thread[(739*4)+1] <= 1'b1;
                  active_thread[(739*4)+2] <= 1'b1;
                  active_thread[(739*4)+3] <= 1'b1;
                  spc739_inst_done         <= `ARIANE_CORE739.piton_pc_vld;
                  spc739_phy_pc_w          <= `ARIANE_CORE739.piton_pc;
                end
            end
    

            assign spc740_thread_id = 2'b00;
            assign spc740_rtl_pc = spc740_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(740*4)]   <= 1'b0;
                  active_thread[(740*4)+1] <= 1'b0;
                  active_thread[(740*4)+2] <= 1'b0;
                  active_thread[(740*4)+3] <= 1'b0;
                  spc740_inst_done         <= 0;
                  spc740_phy_pc_w          <= 0;
                end else begin
                  active_thread[(740*4)]   <= 1'b1;
                  active_thread[(740*4)+1] <= 1'b1;
                  active_thread[(740*4)+2] <= 1'b1;
                  active_thread[(740*4)+3] <= 1'b1;
                  spc740_inst_done         <= `ARIANE_CORE740.piton_pc_vld;
                  spc740_phy_pc_w          <= `ARIANE_CORE740.piton_pc;
                end
            end
    

            assign spc741_thread_id = 2'b00;
            assign spc741_rtl_pc = spc741_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(741*4)]   <= 1'b0;
                  active_thread[(741*4)+1] <= 1'b0;
                  active_thread[(741*4)+2] <= 1'b0;
                  active_thread[(741*4)+3] <= 1'b0;
                  spc741_inst_done         <= 0;
                  spc741_phy_pc_w          <= 0;
                end else begin
                  active_thread[(741*4)]   <= 1'b1;
                  active_thread[(741*4)+1] <= 1'b1;
                  active_thread[(741*4)+2] <= 1'b1;
                  active_thread[(741*4)+3] <= 1'b1;
                  spc741_inst_done         <= `ARIANE_CORE741.piton_pc_vld;
                  spc741_phy_pc_w          <= `ARIANE_CORE741.piton_pc;
                end
            end
    

            assign spc742_thread_id = 2'b00;
            assign spc742_rtl_pc = spc742_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(742*4)]   <= 1'b0;
                  active_thread[(742*4)+1] <= 1'b0;
                  active_thread[(742*4)+2] <= 1'b0;
                  active_thread[(742*4)+3] <= 1'b0;
                  spc742_inst_done         <= 0;
                  spc742_phy_pc_w          <= 0;
                end else begin
                  active_thread[(742*4)]   <= 1'b1;
                  active_thread[(742*4)+1] <= 1'b1;
                  active_thread[(742*4)+2] <= 1'b1;
                  active_thread[(742*4)+3] <= 1'b1;
                  spc742_inst_done         <= `ARIANE_CORE742.piton_pc_vld;
                  spc742_phy_pc_w          <= `ARIANE_CORE742.piton_pc;
                end
            end
    

            assign spc743_thread_id = 2'b00;
            assign spc743_rtl_pc = spc743_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(743*4)]   <= 1'b0;
                  active_thread[(743*4)+1] <= 1'b0;
                  active_thread[(743*4)+2] <= 1'b0;
                  active_thread[(743*4)+3] <= 1'b0;
                  spc743_inst_done         <= 0;
                  spc743_phy_pc_w          <= 0;
                end else begin
                  active_thread[(743*4)]   <= 1'b1;
                  active_thread[(743*4)+1] <= 1'b1;
                  active_thread[(743*4)+2] <= 1'b1;
                  active_thread[(743*4)+3] <= 1'b1;
                  spc743_inst_done         <= `ARIANE_CORE743.piton_pc_vld;
                  spc743_phy_pc_w          <= `ARIANE_CORE743.piton_pc;
                end
            end
    

            assign spc744_thread_id = 2'b00;
            assign spc744_rtl_pc = spc744_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(744*4)]   <= 1'b0;
                  active_thread[(744*4)+1] <= 1'b0;
                  active_thread[(744*4)+2] <= 1'b0;
                  active_thread[(744*4)+3] <= 1'b0;
                  spc744_inst_done         <= 0;
                  spc744_phy_pc_w          <= 0;
                end else begin
                  active_thread[(744*4)]   <= 1'b1;
                  active_thread[(744*4)+1] <= 1'b1;
                  active_thread[(744*4)+2] <= 1'b1;
                  active_thread[(744*4)+3] <= 1'b1;
                  spc744_inst_done         <= `ARIANE_CORE744.piton_pc_vld;
                  spc744_phy_pc_w          <= `ARIANE_CORE744.piton_pc;
                end
            end
    

            assign spc745_thread_id = 2'b00;
            assign spc745_rtl_pc = spc745_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(745*4)]   <= 1'b0;
                  active_thread[(745*4)+1] <= 1'b0;
                  active_thread[(745*4)+2] <= 1'b0;
                  active_thread[(745*4)+3] <= 1'b0;
                  spc745_inst_done         <= 0;
                  spc745_phy_pc_w          <= 0;
                end else begin
                  active_thread[(745*4)]   <= 1'b1;
                  active_thread[(745*4)+1] <= 1'b1;
                  active_thread[(745*4)+2] <= 1'b1;
                  active_thread[(745*4)+3] <= 1'b1;
                  spc745_inst_done         <= `ARIANE_CORE745.piton_pc_vld;
                  spc745_phy_pc_w          <= `ARIANE_CORE745.piton_pc;
                end
            end
    

            assign spc746_thread_id = 2'b00;
            assign spc746_rtl_pc = spc746_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(746*4)]   <= 1'b0;
                  active_thread[(746*4)+1] <= 1'b0;
                  active_thread[(746*4)+2] <= 1'b0;
                  active_thread[(746*4)+3] <= 1'b0;
                  spc746_inst_done         <= 0;
                  spc746_phy_pc_w          <= 0;
                end else begin
                  active_thread[(746*4)]   <= 1'b1;
                  active_thread[(746*4)+1] <= 1'b1;
                  active_thread[(746*4)+2] <= 1'b1;
                  active_thread[(746*4)+3] <= 1'b1;
                  spc746_inst_done         <= `ARIANE_CORE746.piton_pc_vld;
                  spc746_phy_pc_w          <= `ARIANE_CORE746.piton_pc;
                end
            end
    

            assign spc747_thread_id = 2'b00;
            assign spc747_rtl_pc = spc747_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(747*4)]   <= 1'b0;
                  active_thread[(747*4)+1] <= 1'b0;
                  active_thread[(747*4)+2] <= 1'b0;
                  active_thread[(747*4)+3] <= 1'b0;
                  spc747_inst_done         <= 0;
                  spc747_phy_pc_w          <= 0;
                end else begin
                  active_thread[(747*4)]   <= 1'b1;
                  active_thread[(747*4)+1] <= 1'b1;
                  active_thread[(747*4)+2] <= 1'b1;
                  active_thread[(747*4)+3] <= 1'b1;
                  spc747_inst_done         <= `ARIANE_CORE747.piton_pc_vld;
                  spc747_phy_pc_w          <= `ARIANE_CORE747.piton_pc;
                end
            end
    

            assign spc748_thread_id = 2'b00;
            assign spc748_rtl_pc = spc748_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(748*4)]   <= 1'b0;
                  active_thread[(748*4)+1] <= 1'b0;
                  active_thread[(748*4)+2] <= 1'b0;
                  active_thread[(748*4)+3] <= 1'b0;
                  spc748_inst_done         <= 0;
                  spc748_phy_pc_w          <= 0;
                end else begin
                  active_thread[(748*4)]   <= 1'b1;
                  active_thread[(748*4)+1] <= 1'b1;
                  active_thread[(748*4)+2] <= 1'b1;
                  active_thread[(748*4)+3] <= 1'b1;
                  spc748_inst_done         <= `ARIANE_CORE748.piton_pc_vld;
                  spc748_phy_pc_w          <= `ARIANE_CORE748.piton_pc;
                end
            end
    

            assign spc749_thread_id = 2'b00;
            assign spc749_rtl_pc = spc749_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(749*4)]   <= 1'b0;
                  active_thread[(749*4)+1] <= 1'b0;
                  active_thread[(749*4)+2] <= 1'b0;
                  active_thread[(749*4)+3] <= 1'b0;
                  spc749_inst_done         <= 0;
                  spc749_phy_pc_w          <= 0;
                end else begin
                  active_thread[(749*4)]   <= 1'b1;
                  active_thread[(749*4)+1] <= 1'b1;
                  active_thread[(749*4)+2] <= 1'b1;
                  active_thread[(749*4)+3] <= 1'b1;
                  spc749_inst_done         <= `ARIANE_CORE749.piton_pc_vld;
                  spc749_phy_pc_w          <= `ARIANE_CORE749.piton_pc;
                end
            end
    

            assign spc750_thread_id = 2'b00;
            assign spc750_rtl_pc = spc750_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(750*4)]   <= 1'b0;
                  active_thread[(750*4)+1] <= 1'b0;
                  active_thread[(750*4)+2] <= 1'b0;
                  active_thread[(750*4)+3] <= 1'b0;
                  spc750_inst_done         <= 0;
                  spc750_phy_pc_w          <= 0;
                end else begin
                  active_thread[(750*4)]   <= 1'b1;
                  active_thread[(750*4)+1] <= 1'b1;
                  active_thread[(750*4)+2] <= 1'b1;
                  active_thread[(750*4)+3] <= 1'b1;
                  spc750_inst_done         <= `ARIANE_CORE750.piton_pc_vld;
                  spc750_phy_pc_w          <= `ARIANE_CORE750.piton_pc;
                end
            end
    

            assign spc751_thread_id = 2'b00;
            assign spc751_rtl_pc = spc751_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(751*4)]   <= 1'b0;
                  active_thread[(751*4)+1] <= 1'b0;
                  active_thread[(751*4)+2] <= 1'b0;
                  active_thread[(751*4)+3] <= 1'b0;
                  spc751_inst_done         <= 0;
                  spc751_phy_pc_w          <= 0;
                end else begin
                  active_thread[(751*4)]   <= 1'b1;
                  active_thread[(751*4)+1] <= 1'b1;
                  active_thread[(751*4)+2] <= 1'b1;
                  active_thread[(751*4)+3] <= 1'b1;
                  spc751_inst_done         <= `ARIANE_CORE751.piton_pc_vld;
                  spc751_phy_pc_w          <= `ARIANE_CORE751.piton_pc;
                end
            end
    

            assign spc752_thread_id = 2'b00;
            assign spc752_rtl_pc = spc752_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(752*4)]   <= 1'b0;
                  active_thread[(752*4)+1] <= 1'b0;
                  active_thread[(752*4)+2] <= 1'b0;
                  active_thread[(752*4)+3] <= 1'b0;
                  spc752_inst_done         <= 0;
                  spc752_phy_pc_w          <= 0;
                end else begin
                  active_thread[(752*4)]   <= 1'b1;
                  active_thread[(752*4)+1] <= 1'b1;
                  active_thread[(752*4)+2] <= 1'b1;
                  active_thread[(752*4)+3] <= 1'b1;
                  spc752_inst_done         <= `ARIANE_CORE752.piton_pc_vld;
                  spc752_phy_pc_w          <= `ARIANE_CORE752.piton_pc;
                end
            end
    

            assign spc753_thread_id = 2'b00;
            assign spc753_rtl_pc = spc753_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(753*4)]   <= 1'b0;
                  active_thread[(753*4)+1] <= 1'b0;
                  active_thread[(753*4)+2] <= 1'b0;
                  active_thread[(753*4)+3] <= 1'b0;
                  spc753_inst_done         <= 0;
                  spc753_phy_pc_w          <= 0;
                end else begin
                  active_thread[(753*4)]   <= 1'b1;
                  active_thread[(753*4)+1] <= 1'b1;
                  active_thread[(753*4)+2] <= 1'b1;
                  active_thread[(753*4)+3] <= 1'b1;
                  spc753_inst_done         <= `ARIANE_CORE753.piton_pc_vld;
                  spc753_phy_pc_w          <= `ARIANE_CORE753.piton_pc;
                end
            end
    

            assign spc754_thread_id = 2'b00;
            assign spc754_rtl_pc = spc754_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(754*4)]   <= 1'b0;
                  active_thread[(754*4)+1] <= 1'b0;
                  active_thread[(754*4)+2] <= 1'b0;
                  active_thread[(754*4)+3] <= 1'b0;
                  spc754_inst_done         <= 0;
                  spc754_phy_pc_w          <= 0;
                end else begin
                  active_thread[(754*4)]   <= 1'b1;
                  active_thread[(754*4)+1] <= 1'b1;
                  active_thread[(754*4)+2] <= 1'b1;
                  active_thread[(754*4)+3] <= 1'b1;
                  spc754_inst_done         <= `ARIANE_CORE754.piton_pc_vld;
                  spc754_phy_pc_w          <= `ARIANE_CORE754.piton_pc;
                end
            end
    

            assign spc755_thread_id = 2'b00;
            assign spc755_rtl_pc = spc755_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(755*4)]   <= 1'b0;
                  active_thread[(755*4)+1] <= 1'b0;
                  active_thread[(755*4)+2] <= 1'b0;
                  active_thread[(755*4)+3] <= 1'b0;
                  spc755_inst_done         <= 0;
                  spc755_phy_pc_w          <= 0;
                end else begin
                  active_thread[(755*4)]   <= 1'b1;
                  active_thread[(755*4)+1] <= 1'b1;
                  active_thread[(755*4)+2] <= 1'b1;
                  active_thread[(755*4)+3] <= 1'b1;
                  spc755_inst_done         <= `ARIANE_CORE755.piton_pc_vld;
                  spc755_phy_pc_w          <= `ARIANE_CORE755.piton_pc;
                end
            end
    

            assign spc756_thread_id = 2'b00;
            assign spc756_rtl_pc = spc756_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(756*4)]   <= 1'b0;
                  active_thread[(756*4)+1] <= 1'b0;
                  active_thread[(756*4)+2] <= 1'b0;
                  active_thread[(756*4)+3] <= 1'b0;
                  spc756_inst_done         <= 0;
                  spc756_phy_pc_w          <= 0;
                end else begin
                  active_thread[(756*4)]   <= 1'b1;
                  active_thread[(756*4)+1] <= 1'b1;
                  active_thread[(756*4)+2] <= 1'b1;
                  active_thread[(756*4)+3] <= 1'b1;
                  spc756_inst_done         <= `ARIANE_CORE756.piton_pc_vld;
                  spc756_phy_pc_w          <= `ARIANE_CORE756.piton_pc;
                end
            end
    

            assign spc757_thread_id = 2'b00;
            assign spc757_rtl_pc = spc757_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(757*4)]   <= 1'b0;
                  active_thread[(757*4)+1] <= 1'b0;
                  active_thread[(757*4)+2] <= 1'b0;
                  active_thread[(757*4)+3] <= 1'b0;
                  spc757_inst_done         <= 0;
                  spc757_phy_pc_w          <= 0;
                end else begin
                  active_thread[(757*4)]   <= 1'b1;
                  active_thread[(757*4)+1] <= 1'b1;
                  active_thread[(757*4)+2] <= 1'b1;
                  active_thread[(757*4)+3] <= 1'b1;
                  spc757_inst_done         <= `ARIANE_CORE757.piton_pc_vld;
                  spc757_phy_pc_w          <= `ARIANE_CORE757.piton_pc;
                end
            end
    

            assign spc758_thread_id = 2'b00;
            assign spc758_rtl_pc = spc758_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(758*4)]   <= 1'b0;
                  active_thread[(758*4)+1] <= 1'b0;
                  active_thread[(758*4)+2] <= 1'b0;
                  active_thread[(758*4)+3] <= 1'b0;
                  spc758_inst_done         <= 0;
                  spc758_phy_pc_w          <= 0;
                end else begin
                  active_thread[(758*4)]   <= 1'b1;
                  active_thread[(758*4)+1] <= 1'b1;
                  active_thread[(758*4)+2] <= 1'b1;
                  active_thread[(758*4)+3] <= 1'b1;
                  spc758_inst_done         <= `ARIANE_CORE758.piton_pc_vld;
                  spc758_phy_pc_w          <= `ARIANE_CORE758.piton_pc;
                end
            end
    

            assign spc759_thread_id = 2'b00;
            assign spc759_rtl_pc = spc759_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(759*4)]   <= 1'b0;
                  active_thread[(759*4)+1] <= 1'b0;
                  active_thread[(759*4)+2] <= 1'b0;
                  active_thread[(759*4)+3] <= 1'b0;
                  spc759_inst_done         <= 0;
                  spc759_phy_pc_w          <= 0;
                end else begin
                  active_thread[(759*4)]   <= 1'b1;
                  active_thread[(759*4)+1] <= 1'b1;
                  active_thread[(759*4)+2] <= 1'b1;
                  active_thread[(759*4)+3] <= 1'b1;
                  spc759_inst_done         <= `ARIANE_CORE759.piton_pc_vld;
                  spc759_phy_pc_w          <= `ARIANE_CORE759.piton_pc;
                end
            end
    

            assign spc760_thread_id = 2'b00;
            assign spc760_rtl_pc = spc760_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(760*4)]   <= 1'b0;
                  active_thread[(760*4)+1] <= 1'b0;
                  active_thread[(760*4)+2] <= 1'b0;
                  active_thread[(760*4)+3] <= 1'b0;
                  spc760_inst_done         <= 0;
                  spc760_phy_pc_w          <= 0;
                end else begin
                  active_thread[(760*4)]   <= 1'b1;
                  active_thread[(760*4)+1] <= 1'b1;
                  active_thread[(760*4)+2] <= 1'b1;
                  active_thread[(760*4)+3] <= 1'b1;
                  spc760_inst_done         <= `ARIANE_CORE760.piton_pc_vld;
                  spc760_phy_pc_w          <= `ARIANE_CORE760.piton_pc;
                end
            end
    

            assign spc761_thread_id = 2'b00;
            assign spc761_rtl_pc = spc761_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(761*4)]   <= 1'b0;
                  active_thread[(761*4)+1] <= 1'b0;
                  active_thread[(761*4)+2] <= 1'b0;
                  active_thread[(761*4)+3] <= 1'b0;
                  spc761_inst_done         <= 0;
                  spc761_phy_pc_w          <= 0;
                end else begin
                  active_thread[(761*4)]   <= 1'b1;
                  active_thread[(761*4)+1] <= 1'b1;
                  active_thread[(761*4)+2] <= 1'b1;
                  active_thread[(761*4)+3] <= 1'b1;
                  spc761_inst_done         <= `ARIANE_CORE761.piton_pc_vld;
                  spc761_phy_pc_w          <= `ARIANE_CORE761.piton_pc;
                end
            end
    

            assign spc762_thread_id = 2'b00;
            assign spc762_rtl_pc = spc762_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(762*4)]   <= 1'b0;
                  active_thread[(762*4)+1] <= 1'b0;
                  active_thread[(762*4)+2] <= 1'b0;
                  active_thread[(762*4)+3] <= 1'b0;
                  spc762_inst_done         <= 0;
                  spc762_phy_pc_w          <= 0;
                end else begin
                  active_thread[(762*4)]   <= 1'b1;
                  active_thread[(762*4)+1] <= 1'b1;
                  active_thread[(762*4)+2] <= 1'b1;
                  active_thread[(762*4)+3] <= 1'b1;
                  spc762_inst_done         <= `ARIANE_CORE762.piton_pc_vld;
                  spc762_phy_pc_w          <= `ARIANE_CORE762.piton_pc;
                end
            end
    

            assign spc763_thread_id = 2'b00;
            assign spc763_rtl_pc = spc763_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(763*4)]   <= 1'b0;
                  active_thread[(763*4)+1] <= 1'b0;
                  active_thread[(763*4)+2] <= 1'b0;
                  active_thread[(763*4)+3] <= 1'b0;
                  spc763_inst_done         <= 0;
                  spc763_phy_pc_w          <= 0;
                end else begin
                  active_thread[(763*4)]   <= 1'b1;
                  active_thread[(763*4)+1] <= 1'b1;
                  active_thread[(763*4)+2] <= 1'b1;
                  active_thread[(763*4)+3] <= 1'b1;
                  spc763_inst_done         <= `ARIANE_CORE763.piton_pc_vld;
                  spc763_phy_pc_w          <= `ARIANE_CORE763.piton_pc;
                end
            end
    

            assign spc764_thread_id = 2'b00;
            assign spc764_rtl_pc = spc764_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(764*4)]   <= 1'b0;
                  active_thread[(764*4)+1] <= 1'b0;
                  active_thread[(764*4)+2] <= 1'b0;
                  active_thread[(764*4)+3] <= 1'b0;
                  spc764_inst_done         <= 0;
                  spc764_phy_pc_w          <= 0;
                end else begin
                  active_thread[(764*4)]   <= 1'b1;
                  active_thread[(764*4)+1] <= 1'b1;
                  active_thread[(764*4)+2] <= 1'b1;
                  active_thread[(764*4)+3] <= 1'b1;
                  spc764_inst_done         <= `ARIANE_CORE764.piton_pc_vld;
                  spc764_phy_pc_w          <= `ARIANE_CORE764.piton_pc;
                end
            end
    

            assign spc765_thread_id = 2'b00;
            assign spc765_rtl_pc = spc765_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(765*4)]   <= 1'b0;
                  active_thread[(765*4)+1] <= 1'b0;
                  active_thread[(765*4)+2] <= 1'b0;
                  active_thread[(765*4)+3] <= 1'b0;
                  spc765_inst_done         <= 0;
                  spc765_phy_pc_w          <= 0;
                end else begin
                  active_thread[(765*4)]   <= 1'b1;
                  active_thread[(765*4)+1] <= 1'b1;
                  active_thread[(765*4)+2] <= 1'b1;
                  active_thread[(765*4)+3] <= 1'b1;
                  spc765_inst_done         <= `ARIANE_CORE765.piton_pc_vld;
                  spc765_phy_pc_w          <= `ARIANE_CORE765.piton_pc;
                end
            end
    

            assign spc766_thread_id = 2'b00;
            assign spc766_rtl_pc = spc766_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(766*4)]   <= 1'b0;
                  active_thread[(766*4)+1] <= 1'b0;
                  active_thread[(766*4)+2] <= 1'b0;
                  active_thread[(766*4)+3] <= 1'b0;
                  spc766_inst_done         <= 0;
                  spc766_phy_pc_w          <= 0;
                end else begin
                  active_thread[(766*4)]   <= 1'b1;
                  active_thread[(766*4)+1] <= 1'b1;
                  active_thread[(766*4)+2] <= 1'b1;
                  active_thread[(766*4)+3] <= 1'b1;
                  spc766_inst_done         <= `ARIANE_CORE766.piton_pc_vld;
                  spc766_phy_pc_w          <= `ARIANE_CORE766.piton_pc;
                end
            end
    

            assign spc767_thread_id = 2'b00;
            assign spc767_rtl_pc = spc767_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(767*4)]   <= 1'b0;
                  active_thread[(767*4)+1] <= 1'b0;
                  active_thread[(767*4)+2] <= 1'b0;
                  active_thread[(767*4)+3] <= 1'b0;
                  spc767_inst_done         <= 0;
                  spc767_phy_pc_w          <= 0;
                end else begin
                  active_thread[(767*4)]   <= 1'b1;
                  active_thread[(767*4)+1] <= 1'b1;
                  active_thread[(767*4)+2] <= 1'b1;
                  active_thread[(767*4)+3] <= 1'b1;
                  spc767_inst_done         <= `ARIANE_CORE767.piton_pc_vld;
                  spc767_phy_pc_w          <= `ARIANE_CORE767.piton_pc;
                end
            end
    

            assign spc768_thread_id = 2'b00;
            assign spc768_rtl_pc = spc768_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(768*4)]   <= 1'b0;
                  active_thread[(768*4)+1] <= 1'b0;
                  active_thread[(768*4)+2] <= 1'b0;
                  active_thread[(768*4)+3] <= 1'b0;
                  spc768_inst_done         <= 0;
                  spc768_phy_pc_w          <= 0;
                end else begin
                  active_thread[(768*4)]   <= 1'b1;
                  active_thread[(768*4)+1] <= 1'b1;
                  active_thread[(768*4)+2] <= 1'b1;
                  active_thread[(768*4)+3] <= 1'b1;
                  spc768_inst_done         <= `ARIANE_CORE768.piton_pc_vld;
                  spc768_phy_pc_w          <= `ARIANE_CORE768.piton_pc;
                end
            end
    

            assign spc769_thread_id = 2'b00;
            assign spc769_rtl_pc = spc769_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(769*4)]   <= 1'b0;
                  active_thread[(769*4)+1] <= 1'b0;
                  active_thread[(769*4)+2] <= 1'b0;
                  active_thread[(769*4)+3] <= 1'b0;
                  spc769_inst_done         <= 0;
                  spc769_phy_pc_w          <= 0;
                end else begin
                  active_thread[(769*4)]   <= 1'b1;
                  active_thread[(769*4)+1] <= 1'b1;
                  active_thread[(769*4)+2] <= 1'b1;
                  active_thread[(769*4)+3] <= 1'b1;
                  spc769_inst_done         <= `ARIANE_CORE769.piton_pc_vld;
                  spc769_phy_pc_w          <= `ARIANE_CORE769.piton_pc;
                end
            end
    

            assign spc770_thread_id = 2'b00;
            assign spc770_rtl_pc = spc770_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(770*4)]   <= 1'b0;
                  active_thread[(770*4)+1] <= 1'b0;
                  active_thread[(770*4)+2] <= 1'b0;
                  active_thread[(770*4)+3] <= 1'b0;
                  spc770_inst_done         <= 0;
                  spc770_phy_pc_w          <= 0;
                end else begin
                  active_thread[(770*4)]   <= 1'b1;
                  active_thread[(770*4)+1] <= 1'b1;
                  active_thread[(770*4)+2] <= 1'b1;
                  active_thread[(770*4)+3] <= 1'b1;
                  spc770_inst_done         <= `ARIANE_CORE770.piton_pc_vld;
                  spc770_phy_pc_w          <= `ARIANE_CORE770.piton_pc;
                end
            end
    

            assign spc771_thread_id = 2'b00;
            assign spc771_rtl_pc = spc771_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(771*4)]   <= 1'b0;
                  active_thread[(771*4)+1] <= 1'b0;
                  active_thread[(771*4)+2] <= 1'b0;
                  active_thread[(771*4)+3] <= 1'b0;
                  spc771_inst_done         <= 0;
                  spc771_phy_pc_w          <= 0;
                end else begin
                  active_thread[(771*4)]   <= 1'b1;
                  active_thread[(771*4)+1] <= 1'b1;
                  active_thread[(771*4)+2] <= 1'b1;
                  active_thread[(771*4)+3] <= 1'b1;
                  spc771_inst_done         <= `ARIANE_CORE771.piton_pc_vld;
                  spc771_phy_pc_w          <= `ARIANE_CORE771.piton_pc;
                end
            end
    

            assign spc772_thread_id = 2'b00;
            assign spc772_rtl_pc = spc772_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(772*4)]   <= 1'b0;
                  active_thread[(772*4)+1] <= 1'b0;
                  active_thread[(772*4)+2] <= 1'b0;
                  active_thread[(772*4)+3] <= 1'b0;
                  spc772_inst_done         <= 0;
                  spc772_phy_pc_w          <= 0;
                end else begin
                  active_thread[(772*4)]   <= 1'b1;
                  active_thread[(772*4)+1] <= 1'b1;
                  active_thread[(772*4)+2] <= 1'b1;
                  active_thread[(772*4)+3] <= 1'b1;
                  spc772_inst_done         <= `ARIANE_CORE772.piton_pc_vld;
                  spc772_phy_pc_w          <= `ARIANE_CORE772.piton_pc;
                end
            end
    

            assign spc773_thread_id = 2'b00;
            assign spc773_rtl_pc = spc773_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(773*4)]   <= 1'b0;
                  active_thread[(773*4)+1] <= 1'b0;
                  active_thread[(773*4)+2] <= 1'b0;
                  active_thread[(773*4)+3] <= 1'b0;
                  spc773_inst_done         <= 0;
                  spc773_phy_pc_w          <= 0;
                end else begin
                  active_thread[(773*4)]   <= 1'b1;
                  active_thread[(773*4)+1] <= 1'b1;
                  active_thread[(773*4)+2] <= 1'b1;
                  active_thread[(773*4)+3] <= 1'b1;
                  spc773_inst_done         <= `ARIANE_CORE773.piton_pc_vld;
                  spc773_phy_pc_w          <= `ARIANE_CORE773.piton_pc;
                end
            end
    

            assign spc774_thread_id = 2'b00;
            assign spc774_rtl_pc = spc774_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(774*4)]   <= 1'b0;
                  active_thread[(774*4)+1] <= 1'b0;
                  active_thread[(774*4)+2] <= 1'b0;
                  active_thread[(774*4)+3] <= 1'b0;
                  spc774_inst_done         <= 0;
                  spc774_phy_pc_w          <= 0;
                end else begin
                  active_thread[(774*4)]   <= 1'b1;
                  active_thread[(774*4)+1] <= 1'b1;
                  active_thread[(774*4)+2] <= 1'b1;
                  active_thread[(774*4)+3] <= 1'b1;
                  spc774_inst_done         <= `ARIANE_CORE774.piton_pc_vld;
                  spc774_phy_pc_w          <= `ARIANE_CORE774.piton_pc;
                end
            end
    

            assign spc775_thread_id = 2'b00;
            assign spc775_rtl_pc = spc775_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(775*4)]   <= 1'b0;
                  active_thread[(775*4)+1] <= 1'b0;
                  active_thread[(775*4)+2] <= 1'b0;
                  active_thread[(775*4)+3] <= 1'b0;
                  spc775_inst_done         <= 0;
                  spc775_phy_pc_w          <= 0;
                end else begin
                  active_thread[(775*4)]   <= 1'b1;
                  active_thread[(775*4)+1] <= 1'b1;
                  active_thread[(775*4)+2] <= 1'b1;
                  active_thread[(775*4)+3] <= 1'b1;
                  spc775_inst_done         <= `ARIANE_CORE775.piton_pc_vld;
                  spc775_phy_pc_w          <= `ARIANE_CORE775.piton_pc;
                end
            end
    

            assign spc776_thread_id = 2'b00;
            assign spc776_rtl_pc = spc776_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(776*4)]   <= 1'b0;
                  active_thread[(776*4)+1] <= 1'b0;
                  active_thread[(776*4)+2] <= 1'b0;
                  active_thread[(776*4)+3] <= 1'b0;
                  spc776_inst_done         <= 0;
                  spc776_phy_pc_w          <= 0;
                end else begin
                  active_thread[(776*4)]   <= 1'b1;
                  active_thread[(776*4)+1] <= 1'b1;
                  active_thread[(776*4)+2] <= 1'b1;
                  active_thread[(776*4)+3] <= 1'b1;
                  spc776_inst_done         <= `ARIANE_CORE776.piton_pc_vld;
                  spc776_phy_pc_w          <= `ARIANE_CORE776.piton_pc;
                end
            end
    

            assign spc777_thread_id = 2'b00;
            assign spc777_rtl_pc = spc777_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(777*4)]   <= 1'b0;
                  active_thread[(777*4)+1] <= 1'b0;
                  active_thread[(777*4)+2] <= 1'b0;
                  active_thread[(777*4)+3] <= 1'b0;
                  spc777_inst_done         <= 0;
                  spc777_phy_pc_w          <= 0;
                end else begin
                  active_thread[(777*4)]   <= 1'b1;
                  active_thread[(777*4)+1] <= 1'b1;
                  active_thread[(777*4)+2] <= 1'b1;
                  active_thread[(777*4)+3] <= 1'b1;
                  spc777_inst_done         <= `ARIANE_CORE777.piton_pc_vld;
                  spc777_phy_pc_w          <= `ARIANE_CORE777.piton_pc;
                end
            end
    

            assign spc778_thread_id = 2'b00;
            assign spc778_rtl_pc = spc778_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(778*4)]   <= 1'b0;
                  active_thread[(778*4)+1] <= 1'b0;
                  active_thread[(778*4)+2] <= 1'b0;
                  active_thread[(778*4)+3] <= 1'b0;
                  spc778_inst_done         <= 0;
                  spc778_phy_pc_w          <= 0;
                end else begin
                  active_thread[(778*4)]   <= 1'b1;
                  active_thread[(778*4)+1] <= 1'b1;
                  active_thread[(778*4)+2] <= 1'b1;
                  active_thread[(778*4)+3] <= 1'b1;
                  spc778_inst_done         <= `ARIANE_CORE778.piton_pc_vld;
                  spc778_phy_pc_w          <= `ARIANE_CORE778.piton_pc;
                end
            end
    

            assign spc779_thread_id = 2'b00;
            assign spc779_rtl_pc = spc779_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(779*4)]   <= 1'b0;
                  active_thread[(779*4)+1] <= 1'b0;
                  active_thread[(779*4)+2] <= 1'b0;
                  active_thread[(779*4)+3] <= 1'b0;
                  spc779_inst_done         <= 0;
                  spc779_phy_pc_w          <= 0;
                end else begin
                  active_thread[(779*4)]   <= 1'b1;
                  active_thread[(779*4)+1] <= 1'b1;
                  active_thread[(779*4)+2] <= 1'b1;
                  active_thread[(779*4)+3] <= 1'b1;
                  spc779_inst_done         <= `ARIANE_CORE779.piton_pc_vld;
                  spc779_phy_pc_w          <= `ARIANE_CORE779.piton_pc;
                end
            end
    

            assign spc780_thread_id = 2'b00;
            assign spc780_rtl_pc = spc780_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(780*4)]   <= 1'b0;
                  active_thread[(780*4)+1] <= 1'b0;
                  active_thread[(780*4)+2] <= 1'b0;
                  active_thread[(780*4)+3] <= 1'b0;
                  spc780_inst_done         <= 0;
                  spc780_phy_pc_w          <= 0;
                end else begin
                  active_thread[(780*4)]   <= 1'b1;
                  active_thread[(780*4)+1] <= 1'b1;
                  active_thread[(780*4)+2] <= 1'b1;
                  active_thread[(780*4)+3] <= 1'b1;
                  spc780_inst_done         <= `ARIANE_CORE780.piton_pc_vld;
                  spc780_phy_pc_w          <= `ARIANE_CORE780.piton_pc;
                end
            end
    

            assign spc781_thread_id = 2'b00;
            assign spc781_rtl_pc = spc781_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(781*4)]   <= 1'b0;
                  active_thread[(781*4)+1] <= 1'b0;
                  active_thread[(781*4)+2] <= 1'b0;
                  active_thread[(781*4)+3] <= 1'b0;
                  spc781_inst_done         <= 0;
                  spc781_phy_pc_w          <= 0;
                end else begin
                  active_thread[(781*4)]   <= 1'b1;
                  active_thread[(781*4)+1] <= 1'b1;
                  active_thread[(781*4)+2] <= 1'b1;
                  active_thread[(781*4)+3] <= 1'b1;
                  spc781_inst_done         <= `ARIANE_CORE781.piton_pc_vld;
                  spc781_phy_pc_w          <= `ARIANE_CORE781.piton_pc;
                end
            end
    

            assign spc782_thread_id = 2'b00;
            assign spc782_rtl_pc = spc782_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(782*4)]   <= 1'b0;
                  active_thread[(782*4)+1] <= 1'b0;
                  active_thread[(782*4)+2] <= 1'b0;
                  active_thread[(782*4)+3] <= 1'b0;
                  spc782_inst_done         <= 0;
                  spc782_phy_pc_w          <= 0;
                end else begin
                  active_thread[(782*4)]   <= 1'b1;
                  active_thread[(782*4)+1] <= 1'b1;
                  active_thread[(782*4)+2] <= 1'b1;
                  active_thread[(782*4)+3] <= 1'b1;
                  spc782_inst_done         <= `ARIANE_CORE782.piton_pc_vld;
                  spc782_phy_pc_w          <= `ARIANE_CORE782.piton_pc;
                end
            end
    

            assign spc783_thread_id = 2'b00;
            assign spc783_rtl_pc = spc783_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(783*4)]   <= 1'b0;
                  active_thread[(783*4)+1] <= 1'b0;
                  active_thread[(783*4)+2] <= 1'b0;
                  active_thread[(783*4)+3] <= 1'b0;
                  spc783_inst_done         <= 0;
                  spc783_phy_pc_w          <= 0;
                end else begin
                  active_thread[(783*4)]   <= 1'b1;
                  active_thread[(783*4)+1] <= 1'b1;
                  active_thread[(783*4)+2] <= 1'b1;
                  active_thread[(783*4)+3] <= 1'b1;
                  spc783_inst_done         <= `ARIANE_CORE783.piton_pc_vld;
                  spc783_phy_pc_w          <= `ARIANE_CORE783.piton_pc;
                end
            end
    

            assign spc784_thread_id = 2'b00;
            assign spc784_rtl_pc = spc784_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(784*4)]   <= 1'b0;
                  active_thread[(784*4)+1] <= 1'b0;
                  active_thread[(784*4)+2] <= 1'b0;
                  active_thread[(784*4)+3] <= 1'b0;
                  spc784_inst_done         <= 0;
                  spc784_phy_pc_w          <= 0;
                end else begin
                  active_thread[(784*4)]   <= 1'b1;
                  active_thread[(784*4)+1] <= 1'b1;
                  active_thread[(784*4)+2] <= 1'b1;
                  active_thread[(784*4)+3] <= 1'b1;
                  spc784_inst_done         <= `ARIANE_CORE784.piton_pc_vld;
                  spc784_phy_pc_w          <= `ARIANE_CORE784.piton_pc;
                end
            end
    

            assign spc785_thread_id = 2'b00;
            assign spc785_rtl_pc = spc785_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(785*4)]   <= 1'b0;
                  active_thread[(785*4)+1] <= 1'b0;
                  active_thread[(785*4)+2] <= 1'b0;
                  active_thread[(785*4)+3] <= 1'b0;
                  spc785_inst_done         <= 0;
                  spc785_phy_pc_w          <= 0;
                end else begin
                  active_thread[(785*4)]   <= 1'b1;
                  active_thread[(785*4)+1] <= 1'b1;
                  active_thread[(785*4)+2] <= 1'b1;
                  active_thread[(785*4)+3] <= 1'b1;
                  spc785_inst_done         <= `ARIANE_CORE785.piton_pc_vld;
                  spc785_phy_pc_w          <= `ARIANE_CORE785.piton_pc;
                end
            end
    

            assign spc786_thread_id = 2'b00;
            assign spc786_rtl_pc = spc786_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(786*4)]   <= 1'b0;
                  active_thread[(786*4)+1] <= 1'b0;
                  active_thread[(786*4)+2] <= 1'b0;
                  active_thread[(786*4)+3] <= 1'b0;
                  spc786_inst_done         <= 0;
                  spc786_phy_pc_w          <= 0;
                end else begin
                  active_thread[(786*4)]   <= 1'b1;
                  active_thread[(786*4)+1] <= 1'b1;
                  active_thread[(786*4)+2] <= 1'b1;
                  active_thread[(786*4)+3] <= 1'b1;
                  spc786_inst_done         <= `ARIANE_CORE786.piton_pc_vld;
                  spc786_phy_pc_w          <= `ARIANE_CORE786.piton_pc;
                end
            end
    

            assign spc787_thread_id = 2'b00;
            assign spc787_rtl_pc = spc787_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(787*4)]   <= 1'b0;
                  active_thread[(787*4)+1] <= 1'b0;
                  active_thread[(787*4)+2] <= 1'b0;
                  active_thread[(787*4)+3] <= 1'b0;
                  spc787_inst_done         <= 0;
                  spc787_phy_pc_w          <= 0;
                end else begin
                  active_thread[(787*4)]   <= 1'b1;
                  active_thread[(787*4)+1] <= 1'b1;
                  active_thread[(787*4)+2] <= 1'b1;
                  active_thread[(787*4)+3] <= 1'b1;
                  spc787_inst_done         <= `ARIANE_CORE787.piton_pc_vld;
                  spc787_phy_pc_w          <= `ARIANE_CORE787.piton_pc;
                end
            end
    

            assign spc788_thread_id = 2'b00;
            assign spc788_rtl_pc = spc788_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(788*4)]   <= 1'b0;
                  active_thread[(788*4)+1] <= 1'b0;
                  active_thread[(788*4)+2] <= 1'b0;
                  active_thread[(788*4)+3] <= 1'b0;
                  spc788_inst_done         <= 0;
                  spc788_phy_pc_w          <= 0;
                end else begin
                  active_thread[(788*4)]   <= 1'b1;
                  active_thread[(788*4)+1] <= 1'b1;
                  active_thread[(788*4)+2] <= 1'b1;
                  active_thread[(788*4)+3] <= 1'b1;
                  spc788_inst_done         <= `ARIANE_CORE788.piton_pc_vld;
                  spc788_phy_pc_w          <= `ARIANE_CORE788.piton_pc;
                end
            end
    

            assign spc789_thread_id = 2'b00;
            assign spc789_rtl_pc = spc789_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(789*4)]   <= 1'b0;
                  active_thread[(789*4)+1] <= 1'b0;
                  active_thread[(789*4)+2] <= 1'b0;
                  active_thread[(789*4)+3] <= 1'b0;
                  spc789_inst_done         <= 0;
                  spc789_phy_pc_w          <= 0;
                end else begin
                  active_thread[(789*4)]   <= 1'b1;
                  active_thread[(789*4)+1] <= 1'b1;
                  active_thread[(789*4)+2] <= 1'b1;
                  active_thread[(789*4)+3] <= 1'b1;
                  spc789_inst_done         <= `ARIANE_CORE789.piton_pc_vld;
                  spc789_phy_pc_w          <= `ARIANE_CORE789.piton_pc;
                end
            end
    

            assign spc790_thread_id = 2'b00;
            assign spc790_rtl_pc = spc790_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(790*4)]   <= 1'b0;
                  active_thread[(790*4)+1] <= 1'b0;
                  active_thread[(790*4)+2] <= 1'b0;
                  active_thread[(790*4)+3] <= 1'b0;
                  spc790_inst_done         <= 0;
                  spc790_phy_pc_w          <= 0;
                end else begin
                  active_thread[(790*4)]   <= 1'b1;
                  active_thread[(790*4)+1] <= 1'b1;
                  active_thread[(790*4)+2] <= 1'b1;
                  active_thread[(790*4)+3] <= 1'b1;
                  spc790_inst_done         <= `ARIANE_CORE790.piton_pc_vld;
                  spc790_phy_pc_w          <= `ARIANE_CORE790.piton_pc;
                end
            end
    

            assign spc791_thread_id = 2'b00;
            assign spc791_rtl_pc = spc791_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(791*4)]   <= 1'b0;
                  active_thread[(791*4)+1] <= 1'b0;
                  active_thread[(791*4)+2] <= 1'b0;
                  active_thread[(791*4)+3] <= 1'b0;
                  spc791_inst_done         <= 0;
                  spc791_phy_pc_w          <= 0;
                end else begin
                  active_thread[(791*4)]   <= 1'b1;
                  active_thread[(791*4)+1] <= 1'b1;
                  active_thread[(791*4)+2] <= 1'b1;
                  active_thread[(791*4)+3] <= 1'b1;
                  spc791_inst_done         <= `ARIANE_CORE791.piton_pc_vld;
                  spc791_phy_pc_w          <= `ARIANE_CORE791.piton_pc;
                end
            end
    

            assign spc792_thread_id = 2'b00;
            assign spc792_rtl_pc = spc792_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(792*4)]   <= 1'b0;
                  active_thread[(792*4)+1] <= 1'b0;
                  active_thread[(792*4)+2] <= 1'b0;
                  active_thread[(792*4)+3] <= 1'b0;
                  spc792_inst_done         <= 0;
                  spc792_phy_pc_w          <= 0;
                end else begin
                  active_thread[(792*4)]   <= 1'b1;
                  active_thread[(792*4)+1] <= 1'b1;
                  active_thread[(792*4)+2] <= 1'b1;
                  active_thread[(792*4)+3] <= 1'b1;
                  spc792_inst_done         <= `ARIANE_CORE792.piton_pc_vld;
                  spc792_phy_pc_w          <= `ARIANE_CORE792.piton_pc;
                end
            end
    

            assign spc793_thread_id = 2'b00;
            assign spc793_rtl_pc = spc793_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(793*4)]   <= 1'b0;
                  active_thread[(793*4)+1] <= 1'b0;
                  active_thread[(793*4)+2] <= 1'b0;
                  active_thread[(793*4)+3] <= 1'b0;
                  spc793_inst_done         <= 0;
                  spc793_phy_pc_w          <= 0;
                end else begin
                  active_thread[(793*4)]   <= 1'b1;
                  active_thread[(793*4)+1] <= 1'b1;
                  active_thread[(793*4)+2] <= 1'b1;
                  active_thread[(793*4)+3] <= 1'b1;
                  spc793_inst_done         <= `ARIANE_CORE793.piton_pc_vld;
                  spc793_phy_pc_w          <= `ARIANE_CORE793.piton_pc;
                end
            end
    

            assign spc794_thread_id = 2'b00;
            assign spc794_rtl_pc = spc794_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(794*4)]   <= 1'b0;
                  active_thread[(794*4)+1] <= 1'b0;
                  active_thread[(794*4)+2] <= 1'b0;
                  active_thread[(794*4)+3] <= 1'b0;
                  spc794_inst_done         <= 0;
                  spc794_phy_pc_w          <= 0;
                end else begin
                  active_thread[(794*4)]   <= 1'b1;
                  active_thread[(794*4)+1] <= 1'b1;
                  active_thread[(794*4)+2] <= 1'b1;
                  active_thread[(794*4)+3] <= 1'b1;
                  spc794_inst_done         <= `ARIANE_CORE794.piton_pc_vld;
                  spc794_phy_pc_w          <= `ARIANE_CORE794.piton_pc;
                end
            end
    

            assign spc795_thread_id = 2'b00;
            assign spc795_rtl_pc = spc795_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(795*4)]   <= 1'b0;
                  active_thread[(795*4)+1] <= 1'b0;
                  active_thread[(795*4)+2] <= 1'b0;
                  active_thread[(795*4)+3] <= 1'b0;
                  spc795_inst_done         <= 0;
                  spc795_phy_pc_w          <= 0;
                end else begin
                  active_thread[(795*4)]   <= 1'b1;
                  active_thread[(795*4)+1] <= 1'b1;
                  active_thread[(795*4)+2] <= 1'b1;
                  active_thread[(795*4)+3] <= 1'b1;
                  spc795_inst_done         <= `ARIANE_CORE795.piton_pc_vld;
                  spc795_phy_pc_w          <= `ARIANE_CORE795.piton_pc;
                end
            end
    

            assign spc796_thread_id = 2'b00;
            assign spc796_rtl_pc = spc796_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(796*4)]   <= 1'b0;
                  active_thread[(796*4)+1] <= 1'b0;
                  active_thread[(796*4)+2] <= 1'b0;
                  active_thread[(796*4)+3] <= 1'b0;
                  spc796_inst_done         <= 0;
                  spc796_phy_pc_w          <= 0;
                end else begin
                  active_thread[(796*4)]   <= 1'b1;
                  active_thread[(796*4)+1] <= 1'b1;
                  active_thread[(796*4)+2] <= 1'b1;
                  active_thread[(796*4)+3] <= 1'b1;
                  spc796_inst_done         <= `ARIANE_CORE796.piton_pc_vld;
                  spc796_phy_pc_w          <= `ARIANE_CORE796.piton_pc;
                end
            end
    

            assign spc797_thread_id = 2'b00;
            assign spc797_rtl_pc = spc797_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(797*4)]   <= 1'b0;
                  active_thread[(797*4)+1] <= 1'b0;
                  active_thread[(797*4)+2] <= 1'b0;
                  active_thread[(797*4)+3] <= 1'b0;
                  spc797_inst_done         <= 0;
                  spc797_phy_pc_w          <= 0;
                end else begin
                  active_thread[(797*4)]   <= 1'b1;
                  active_thread[(797*4)+1] <= 1'b1;
                  active_thread[(797*4)+2] <= 1'b1;
                  active_thread[(797*4)+3] <= 1'b1;
                  spc797_inst_done         <= `ARIANE_CORE797.piton_pc_vld;
                  spc797_phy_pc_w          <= `ARIANE_CORE797.piton_pc;
                end
            end
    

            assign spc798_thread_id = 2'b00;
            assign spc798_rtl_pc = spc798_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(798*4)]   <= 1'b0;
                  active_thread[(798*4)+1] <= 1'b0;
                  active_thread[(798*4)+2] <= 1'b0;
                  active_thread[(798*4)+3] <= 1'b0;
                  spc798_inst_done         <= 0;
                  spc798_phy_pc_w          <= 0;
                end else begin
                  active_thread[(798*4)]   <= 1'b1;
                  active_thread[(798*4)+1] <= 1'b1;
                  active_thread[(798*4)+2] <= 1'b1;
                  active_thread[(798*4)+3] <= 1'b1;
                  spc798_inst_done         <= `ARIANE_CORE798.piton_pc_vld;
                  spc798_phy_pc_w          <= `ARIANE_CORE798.piton_pc;
                end
            end
    

            assign spc799_thread_id = 2'b00;
            assign spc799_rtl_pc = spc799_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(799*4)]   <= 1'b0;
                  active_thread[(799*4)+1] <= 1'b0;
                  active_thread[(799*4)+2] <= 1'b0;
                  active_thread[(799*4)+3] <= 1'b0;
                  spc799_inst_done         <= 0;
                  spc799_phy_pc_w          <= 0;
                end else begin
                  active_thread[(799*4)]   <= 1'b1;
                  active_thread[(799*4)+1] <= 1'b1;
                  active_thread[(799*4)+2] <= 1'b1;
                  active_thread[(799*4)+3] <= 1'b1;
                  spc799_inst_done         <= `ARIANE_CORE799.piton_pc_vld;
                  spc799_phy_pc_w          <= `ARIANE_CORE799.piton_pc;
                end
            end
    

            assign spc800_thread_id = 2'b00;
            assign spc800_rtl_pc = spc800_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(800*4)]   <= 1'b0;
                  active_thread[(800*4)+1] <= 1'b0;
                  active_thread[(800*4)+2] <= 1'b0;
                  active_thread[(800*4)+3] <= 1'b0;
                  spc800_inst_done         <= 0;
                  spc800_phy_pc_w          <= 0;
                end else begin
                  active_thread[(800*4)]   <= 1'b1;
                  active_thread[(800*4)+1] <= 1'b1;
                  active_thread[(800*4)+2] <= 1'b1;
                  active_thread[(800*4)+3] <= 1'b1;
                  spc800_inst_done         <= `ARIANE_CORE800.piton_pc_vld;
                  spc800_phy_pc_w          <= `ARIANE_CORE800.piton_pc;
                end
            end
    

            assign spc801_thread_id = 2'b00;
            assign spc801_rtl_pc = spc801_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(801*4)]   <= 1'b0;
                  active_thread[(801*4)+1] <= 1'b0;
                  active_thread[(801*4)+2] <= 1'b0;
                  active_thread[(801*4)+3] <= 1'b0;
                  spc801_inst_done         <= 0;
                  spc801_phy_pc_w          <= 0;
                end else begin
                  active_thread[(801*4)]   <= 1'b1;
                  active_thread[(801*4)+1] <= 1'b1;
                  active_thread[(801*4)+2] <= 1'b1;
                  active_thread[(801*4)+3] <= 1'b1;
                  spc801_inst_done         <= `ARIANE_CORE801.piton_pc_vld;
                  spc801_phy_pc_w          <= `ARIANE_CORE801.piton_pc;
                end
            end
    

            assign spc802_thread_id = 2'b00;
            assign spc802_rtl_pc = spc802_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(802*4)]   <= 1'b0;
                  active_thread[(802*4)+1] <= 1'b0;
                  active_thread[(802*4)+2] <= 1'b0;
                  active_thread[(802*4)+3] <= 1'b0;
                  spc802_inst_done         <= 0;
                  spc802_phy_pc_w          <= 0;
                end else begin
                  active_thread[(802*4)]   <= 1'b1;
                  active_thread[(802*4)+1] <= 1'b1;
                  active_thread[(802*4)+2] <= 1'b1;
                  active_thread[(802*4)+3] <= 1'b1;
                  spc802_inst_done         <= `ARIANE_CORE802.piton_pc_vld;
                  spc802_phy_pc_w          <= `ARIANE_CORE802.piton_pc;
                end
            end
    

            assign spc803_thread_id = 2'b00;
            assign spc803_rtl_pc = spc803_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(803*4)]   <= 1'b0;
                  active_thread[(803*4)+1] <= 1'b0;
                  active_thread[(803*4)+2] <= 1'b0;
                  active_thread[(803*4)+3] <= 1'b0;
                  spc803_inst_done         <= 0;
                  spc803_phy_pc_w          <= 0;
                end else begin
                  active_thread[(803*4)]   <= 1'b1;
                  active_thread[(803*4)+1] <= 1'b1;
                  active_thread[(803*4)+2] <= 1'b1;
                  active_thread[(803*4)+3] <= 1'b1;
                  spc803_inst_done         <= `ARIANE_CORE803.piton_pc_vld;
                  spc803_phy_pc_w          <= `ARIANE_CORE803.piton_pc;
                end
            end
    

            assign spc804_thread_id = 2'b00;
            assign spc804_rtl_pc = spc804_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(804*4)]   <= 1'b0;
                  active_thread[(804*4)+1] <= 1'b0;
                  active_thread[(804*4)+2] <= 1'b0;
                  active_thread[(804*4)+3] <= 1'b0;
                  spc804_inst_done         <= 0;
                  spc804_phy_pc_w          <= 0;
                end else begin
                  active_thread[(804*4)]   <= 1'b1;
                  active_thread[(804*4)+1] <= 1'b1;
                  active_thread[(804*4)+2] <= 1'b1;
                  active_thread[(804*4)+3] <= 1'b1;
                  spc804_inst_done         <= `ARIANE_CORE804.piton_pc_vld;
                  spc804_phy_pc_w          <= `ARIANE_CORE804.piton_pc;
                end
            end
    

            assign spc805_thread_id = 2'b00;
            assign spc805_rtl_pc = spc805_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(805*4)]   <= 1'b0;
                  active_thread[(805*4)+1] <= 1'b0;
                  active_thread[(805*4)+2] <= 1'b0;
                  active_thread[(805*4)+3] <= 1'b0;
                  spc805_inst_done         <= 0;
                  spc805_phy_pc_w          <= 0;
                end else begin
                  active_thread[(805*4)]   <= 1'b1;
                  active_thread[(805*4)+1] <= 1'b1;
                  active_thread[(805*4)+2] <= 1'b1;
                  active_thread[(805*4)+3] <= 1'b1;
                  spc805_inst_done         <= `ARIANE_CORE805.piton_pc_vld;
                  spc805_phy_pc_w          <= `ARIANE_CORE805.piton_pc;
                end
            end
    

            assign spc806_thread_id = 2'b00;
            assign spc806_rtl_pc = spc806_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(806*4)]   <= 1'b0;
                  active_thread[(806*4)+1] <= 1'b0;
                  active_thread[(806*4)+2] <= 1'b0;
                  active_thread[(806*4)+3] <= 1'b0;
                  spc806_inst_done         <= 0;
                  spc806_phy_pc_w          <= 0;
                end else begin
                  active_thread[(806*4)]   <= 1'b1;
                  active_thread[(806*4)+1] <= 1'b1;
                  active_thread[(806*4)+2] <= 1'b1;
                  active_thread[(806*4)+3] <= 1'b1;
                  spc806_inst_done         <= `ARIANE_CORE806.piton_pc_vld;
                  spc806_phy_pc_w          <= `ARIANE_CORE806.piton_pc;
                end
            end
    

            assign spc807_thread_id = 2'b00;
            assign spc807_rtl_pc = spc807_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(807*4)]   <= 1'b0;
                  active_thread[(807*4)+1] <= 1'b0;
                  active_thread[(807*4)+2] <= 1'b0;
                  active_thread[(807*4)+3] <= 1'b0;
                  spc807_inst_done         <= 0;
                  spc807_phy_pc_w          <= 0;
                end else begin
                  active_thread[(807*4)]   <= 1'b1;
                  active_thread[(807*4)+1] <= 1'b1;
                  active_thread[(807*4)+2] <= 1'b1;
                  active_thread[(807*4)+3] <= 1'b1;
                  spc807_inst_done         <= `ARIANE_CORE807.piton_pc_vld;
                  spc807_phy_pc_w          <= `ARIANE_CORE807.piton_pc;
                end
            end
    

            assign spc808_thread_id = 2'b00;
            assign spc808_rtl_pc = spc808_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(808*4)]   <= 1'b0;
                  active_thread[(808*4)+1] <= 1'b0;
                  active_thread[(808*4)+2] <= 1'b0;
                  active_thread[(808*4)+3] <= 1'b0;
                  spc808_inst_done         <= 0;
                  spc808_phy_pc_w          <= 0;
                end else begin
                  active_thread[(808*4)]   <= 1'b1;
                  active_thread[(808*4)+1] <= 1'b1;
                  active_thread[(808*4)+2] <= 1'b1;
                  active_thread[(808*4)+3] <= 1'b1;
                  spc808_inst_done         <= `ARIANE_CORE808.piton_pc_vld;
                  spc808_phy_pc_w          <= `ARIANE_CORE808.piton_pc;
                end
            end
    

            assign spc809_thread_id = 2'b00;
            assign spc809_rtl_pc = spc809_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(809*4)]   <= 1'b0;
                  active_thread[(809*4)+1] <= 1'b0;
                  active_thread[(809*4)+2] <= 1'b0;
                  active_thread[(809*4)+3] <= 1'b0;
                  spc809_inst_done         <= 0;
                  spc809_phy_pc_w          <= 0;
                end else begin
                  active_thread[(809*4)]   <= 1'b1;
                  active_thread[(809*4)+1] <= 1'b1;
                  active_thread[(809*4)+2] <= 1'b1;
                  active_thread[(809*4)+3] <= 1'b1;
                  spc809_inst_done         <= `ARIANE_CORE809.piton_pc_vld;
                  spc809_phy_pc_w          <= `ARIANE_CORE809.piton_pc;
                end
            end
    

            assign spc810_thread_id = 2'b00;
            assign spc810_rtl_pc = spc810_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(810*4)]   <= 1'b0;
                  active_thread[(810*4)+1] <= 1'b0;
                  active_thread[(810*4)+2] <= 1'b0;
                  active_thread[(810*4)+3] <= 1'b0;
                  spc810_inst_done         <= 0;
                  spc810_phy_pc_w          <= 0;
                end else begin
                  active_thread[(810*4)]   <= 1'b1;
                  active_thread[(810*4)+1] <= 1'b1;
                  active_thread[(810*4)+2] <= 1'b1;
                  active_thread[(810*4)+3] <= 1'b1;
                  spc810_inst_done         <= `ARIANE_CORE810.piton_pc_vld;
                  spc810_phy_pc_w          <= `ARIANE_CORE810.piton_pc;
                end
            end
    

            assign spc811_thread_id = 2'b00;
            assign spc811_rtl_pc = spc811_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(811*4)]   <= 1'b0;
                  active_thread[(811*4)+1] <= 1'b0;
                  active_thread[(811*4)+2] <= 1'b0;
                  active_thread[(811*4)+3] <= 1'b0;
                  spc811_inst_done         <= 0;
                  spc811_phy_pc_w          <= 0;
                end else begin
                  active_thread[(811*4)]   <= 1'b1;
                  active_thread[(811*4)+1] <= 1'b1;
                  active_thread[(811*4)+2] <= 1'b1;
                  active_thread[(811*4)+3] <= 1'b1;
                  spc811_inst_done         <= `ARIANE_CORE811.piton_pc_vld;
                  spc811_phy_pc_w          <= `ARIANE_CORE811.piton_pc;
                end
            end
    

            assign spc812_thread_id = 2'b00;
            assign spc812_rtl_pc = spc812_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(812*4)]   <= 1'b0;
                  active_thread[(812*4)+1] <= 1'b0;
                  active_thread[(812*4)+2] <= 1'b0;
                  active_thread[(812*4)+3] <= 1'b0;
                  spc812_inst_done         <= 0;
                  spc812_phy_pc_w          <= 0;
                end else begin
                  active_thread[(812*4)]   <= 1'b1;
                  active_thread[(812*4)+1] <= 1'b1;
                  active_thread[(812*4)+2] <= 1'b1;
                  active_thread[(812*4)+3] <= 1'b1;
                  spc812_inst_done         <= `ARIANE_CORE812.piton_pc_vld;
                  spc812_phy_pc_w          <= `ARIANE_CORE812.piton_pc;
                end
            end
    

            assign spc813_thread_id = 2'b00;
            assign spc813_rtl_pc = spc813_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(813*4)]   <= 1'b0;
                  active_thread[(813*4)+1] <= 1'b0;
                  active_thread[(813*4)+2] <= 1'b0;
                  active_thread[(813*4)+3] <= 1'b0;
                  spc813_inst_done         <= 0;
                  spc813_phy_pc_w          <= 0;
                end else begin
                  active_thread[(813*4)]   <= 1'b1;
                  active_thread[(813*4)+1] <= 1'b1;
                  active_thread[(813*4)+2] <= 1'b1;
                  active_thread[(813*4)+3] <= 1'b1;
                  spc813_inst_done         <= `ARIANE_CORE813.piton_pc_vld;
                  spc813_phy_pc_w          <= `ARIANE_CORE813.piton_pc;
                end
            end
    

            assign spc814_thread_id = 2'b00;
            assign spc814_rtl_pc = spc814_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(814*4)]   <= 1'b0;
                  active_thread[(814*4)+1] <= 1'b0;
                  active_thread[(814*4)+2] <= 1'b0;
                  active_thread[(814*4)+3] <= 1'b0;
                  spc814_inst_done         <= 0;
                  spc814_phy_pc_w          <= 0;
                end else begin
                  active_thread[(814*4)]   <= 1'b1;
                  active_thread[(814*4)+1] <= 1'b1;
                  active_thread[(814*4)+2] <= 1'b1;
                  active_thread[(814*4)+3] <= 1'b1;
                  spc814_inst_done         <= `ARIANE_CORE814.piton_pc_vld;
                  spc814_phy_pc_w          <= `ARIANE_CORE814.piton_pc;
                end
            end
    

            assign spc815_thread_id = 2'b00;
            assign spc815_rtl_pc = spc815_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(815*4)]   <= 1'b0;
                  active_thread[(815*4)+1] <= 1'b0;
                  active_thread[(815*4)+2] <= 1'b0;
                  active_thread[(815*4)+3] <= 1'b0;
                  spc815_inst_done         <= 0;
                  spc815_phy_pc_w          <= 0;
                end else begin
                  active_thread[(815*4)]   <= 1'b1;
                  active_thread[(815*4)+1] <= 1'b1;
                  active_thread[(815*4)+2] <= 1'b1;
                  active_thread[(815*4)+3] <= 1'b1;
                  spc815_inst_done         <= `ARIANE_CORE815.piton_pc_vld;
                  spc815_phy_pc_w          <= `ARIANE_CORE815.piton_pc;
                end
            end
    

            assign spc816_thread_id = 2'b00;
            assign spc816_rtl_pc = spc816_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(816*4)]   <= 1'b0;
                  active_thread[(816*4)+1] <= 1'b0;
                  active_thread[(816*4)+2] <= 1'b0;
                  active_thread[(816*4)+3] <= 1'b0;
                  spc816_inst_done         <= 0;
                  spc816_phy_pc_w          <= 0;
                end else begin
                  active_thread[(816*4)]   <= 1'b1;
                  active_thread[(816*4)+1] <= 1'b1;
                  active_thread[(816*4)+2] <= 1'b1;
                  active_thread[(816*4)+3] <= 1'b1;
                  spc816_inst_done         <= `ARIANE_CORE816.piton_pc_vld;
                  spc816_phy_pc_w          <= `ARIANE_CORE816.piton_pc;
                end
            end
    

            assign spc817_thread_id = 2'b00;
            assign spc817_rtl_pc = spc817_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(817*4)]   <= 1'b0;
                  active_thread[(817*4)+1] <= 1'b0;
                  active_thread[(817*4)+2] <= 1'b0;
                  active_thread[(817*4)+3] <= 1'b0;
                  spc817_inst_done         <= 0;
                  spc817_phy_pc_w          <= 0;
                end else begin
                  active_thread[(817*4)]   <= 1'b1;
                  active_thread[(817*4)+1] <= 1'b1;
                  active_thread[(817*4)+2] <= 1'b1;
                  active_thread[(817*4)+3] <= 1'b1;
                  spc817_inst_done         <= `ARIANE_CORE817.piton_pc_vld;
                  spc817_phy_pc_w          <= `ARIANE_CORE817.piton_pc;
                end
            end
    

            assign spc818_thread_id = 2'b00;
            assign spc818_rtl_pc = spc818_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(818*4)]   <= 1'b0;
                  active_thread[(818*4)+1] <= 1'b0;
                  active_thread[(818*4)+2] <= 1'b0;
                  active_thread[(818*4)+3] <= 1'b0;
                  spc818_inst_done         <= 0;
                  spc818_phy_pc_w          <= 0;
                end else begin
                  active_thread[(818*4)]   <= 1'b1;
                  active_thread[(818*4)+1] <= 1'b1;
                  active_thread[(818*4)+2] <= 1'b1;
                  active_thread[(818*4)+3] <= 1'b1;
                  spc818_inst_done         <= `ARIANE_CORE818.piton_pc_vld;
                  spc818_phy_pc_w          <= `ARIANE_CORE818.piton_pc;
                end
            end
    

            assign spc819_thread_id = 2'b00;
            assign spc819_rtl_pc = spc819_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(819*4)]   <= 1'b0;
                  active_thread[(819*4)+1] <= 1'b0;
                  active_thread[(819*4)+2] <= 1'b0;
                  active_thread[(819*4)+3] <= 1'b0;
                  spc819_inst_done         <= 0;
                  spc819_phy_pc_w          <= 0;
                end else begin
                  active_thread[(819*4)]   <= 1'b1;
                  active_thread[(819*4)+1] <= 1'b1;
                  active_thread[(819*4)+2] <= 1'b1;
                  active_thread[(819*4)+3] <= 1'b1;
                  spc819_inst_done         <= `ARIANE_CORE819.piton_pc_vld;
                  spc819_phy_pc_w          <= `ARIANE_CORE819.piton_pc;
                end
            end
    

            assign spc820_thread_id = 2'b00;
            assign spc820_rtl_pc = spc820_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(820*4)]   <= 1'b0;
                  active_thread[(820*4)+1] <= 1'b0;
                  active_thread[(820*4)+2] <= 1'b0;
                  active_thread[(820*4)+3] <= 1'b0;
                  spc820_inst_done         <= 0;
                  spc820_phy_pc_w          <= 0;
                end else begin
                  active_thread[(820*4)]   <= 1'b1;
                  active_thread[(820*4)+1] <= 1'b1;
                  active_thread[(820*4)+2] <= 1'b1;
                  active_thread[(820*4)+3] <= 1'b1;
                  spc820_inst_done         <= `ARIANE_CORE820.piton_pc_vld;
                  spc820_phy_pc_w          <= `ARIANE_CORE820.piton_pc;
                end
            end
    

            assign spc821_thread_id = 2'b00;
            assign spc821_rtl_pc = spc821_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(821*4)]   <= 1'b0;
                  active_thread[(821*4)+1] <= 1'b0;
                  active_thread[(821*4)+2] <= 1'b0;
                  active_thread[(821*4)+3] <= 1'b0;
                  spc821_inst_done         <= 0;
                  spc821_phy_pc_w          <= 0;
                end else begin
                  active_thread[(821*4)]   <= 1'b1;
                  active_thread[(821*4)+1] <= 1'b1;
                  active_thread[(821*4)+2] <= 1'b1;
                  active_thread[(821*4)+3] <= 1'b1;
                  spc821_inst_done         <= `ARIANE_CORE821.piton_pc_vld;
                  spc821_phy_pc_w          <= `ARIANE_CORE821.piton_pc;
                end
            end
    

            assign spc822_thread_id = 2'b00;
            assign spc822_rtl_pc = spc822_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(822*4)]   <= 1'b0;
                  active_thread[(822*4)+1] <= 1'b0;
                  active_thread[(822*4)+2] <= 1'b0;
                  active_thread[(822*4)+3] <= 1'b0;
                  spc822_inst_done         <= 0;
                  spc822_phy_pc_w          <= 0;
                end else begin
                  active_thread[(822*4)]   <= 1'b1;
                  active_thread[(822*4)+1] <= 1'b1;
                  active_thread[(822*4)+2] <= 1'b1;
                  active_thread[(822*4)+3] <= 1'b1;
                  spc822_inst_done         <= `ARIANE_CORE822.piton_pc_vld;
                  spc822_phy_pc_w          <= `ARIANE_CORE822.piton_pc;
                end
            end
    

            assign spc823_thread_id = 2'b00;
            assign spc823_rtl_pc = spc823_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(823*4)]   <= 1'b0;
                  active_thread[(823*4)+1] <= 1'b0;
                  active_thread[(823*4)+2] <= 1'b0;
                  active_thread[(823*4)+3] <= 1'b0;
                  spc823_inst_done         <= 0;
                  spc823_phy_pc_w          <= 0;
                end else begin
                  active_thread[(823*4)]   <= 1'b1;
                  active_thread[(823*4)+1] <= 1'b1;
                  active_thread[(823*4)+2] <= 1'b1;
                  active_thread[(823*4)+3] <= 1'b1;
                  spc823_inst_done         <= `ARIANE_CORE823.piton_pc_vld;
                  spc823_phy_pc_w          <= `ARIANE_CORE823.piton_pc;
                end
            end
    

            assign spc824_thread_id = 2'b00;
            assign spc824_rtl_pc = spc824_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(824*4)]   <= 1'b0;
                  active_thread[(824*4)+1] <= 1'b0;
                  active_thread[(824*4)+2] <= 1'b0;
                  active_thread[(824*4)+3] <= 1'b0;
                  spc824_inst_done         <= 0;
                  spc824_phy_pc_w          <= 0;
                end else begin
                  active_thread[(824*4)]   <= 1'b1;
                  active_thread[(824*4)+1] <= 1'b1;
                  active_thread[(824*4)+2] <= 1'b1;
                  active_thread[(824*4)+3] <= 1'b1;
                  spc824_inst_done         <= `ARIANE_CORE824.piton_pc_vld;
                  spc824_phy_pc_w          <= `ARIANE_CORE824.piton_pc;
                end
            end
    

            assign spc825_thread_id = 2'b00;
            assign spc825_rtl_pc = spc825_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(825*4)]   <= 1'b0;
                  active_thread[(825*4)+1] <= 1'b0;
                  active_thread[(825*4)+2] <= 1'b0;
                  active_thread[(825*4)+3] <= 1'b0;
                  spc825_inst_done         <= 0;
                  spc825_phy_pc_w          <= 0;
                end else begin
                  active_thread[(825*4)]   <= 1'b1;
                  active_thread[(825*4)+1] <= 1'b1;
                  active_thread[(825*4)+2] <= 1'b1;
                  active_thread[(825*4)+3] <= 1'b1;
                  spc825_inst_done         <= `ARIANE_CORE825.piton_pc_vld;
                  spc825_phy_pc_w          <= `ARIANE_CORE825.piton_pc;
                end
            end
    

            assign spc826_thread_id = 2'b00;
            assign spc826_rtl_pc = spc826_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(826*4)]   <= 1'b0;
                  active_thread[(826*4)+1] <= 1'b0;
                  active_thread[(826*4)+2] <= 1'b0;
                  active_thread[(826*4)+3] <= 1'b0;
                  spc826_inst_done         <= 0;
                  spc826_phy_pc_w          <= 0;
                end else begin
                  active_thread[(826*4)]   <= 1'b1;
                  active_thread[(826*4)+1] <= 1'b1;
                  active_thread[(826*4)+2] <= 1'b1;
                  active_thread[(826*4)+3] <= 1'b1;
                  spc826_inst_done         <= `ARIANE_CORE826.piton_pc_vld;
                  spc826_phy_pc_w          <= `ARIANE_CORE826.piton_pc;
                end
            end
    

            assign spc827_thread_id = 2'b00;
            assign spc827_rtl_pc = spc827_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(827*4)]   <= 1'b0;
                  active_thread[(827*4)+1] <= 1'b0;
                  active_thread[(827*4)+2] <= 1'b0;
                  active_thread[(827*4)+3] <= 1'b0;
                  spc827_inst_done         <= 0;
                  spc827_phy_pc_w          <= 0;
                end else begin
                  active_thread[(827*4)]   <= 1'b1;
                  active_thread[(827*4)+1] <= 1'b1;
                  active_thread[(827*4)+2] <= 1'b1;
                  active_thread[(827*4)+3] <= 1'b1;
                  spc827_inst_done         <= `ARIANE_CORE827.piton_pc_vld;
                  spc827_phy_pc_w          <= `ARIANE_CORE827.piton_pc;
                end
            end
    

            assign spc828_thread_id = 2'b00;
            assign spc828_rtl_pc = spc828_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(828*4)]   <= 1'b0;
                  active_thread[(828*4)+1] <= 1'b0;
                  active_thread[(828*4)+2] <= 1'b0;
                  active_thread[(828*4)+3] <= 1'b0;
                  spc828_inst_done         <= 0;
                  spc828_phy_pc_w          <= 0;
                end else begin
                  active_thread[(828*4)]   <= 1'b1;
                  active_thread[(828*4)+1] <= 1'b1;
                  active_thread[(828*4)+2] <= 1'b1;
                  active_thread[(828*4)+3] <= 1'b1;
                  spc828_inst_done         <= `ARIANE_CORE828.piton_pc_vld;
                  spc828_phy_pc_w          <= `ARIANE_CORE828.piton_pc;
                end
            end
    

            assign spc829_thread_id = 2'b00;
            assign spc829_rtl_pc = spc829_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(829*4)]   <= 1'b0;
                  active_thread[(829*4)+1] <= 1'b0;
                  active_thread[(829*4)+2] <= 1'b0;
                  active_thread[(829*4)+3] <= 1'b0;
                  spc829_inst_done         <= 0;
                  spc829_phy_pc_w          <= 0;
                end else begin
                  active_thread[(829*4)]   <= 1'b1;
                  active_thread[(829*4)+1] <= 1'b1;
                  active_thread[(829*4)+2] <= 1'b1;
                  active_thread[(829*4)+3] <= 1'b1;
                  spc829_inst_done         <= `ARIANE_CORE829.piton_pc_vld;
                  spc829_phy_pc_w          <= `ARIANE_CORE829.piton_pc;
                end
            end
    

            assign spc830_thread_id = 2'b00;
            assign spc830_rtl_pc = spc830_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(830*4)]   <= 1'b0;
                  active_thread[(830*4)+1] <= 1'b0;
                  active_thread[(830*4)+2] <= 1'b0;
                  active_thread[(830*4)+3] <= 1'b0;
                  spc830_inst_done         <= 0;
                  spc830_phy_pc_w          <= 0;
                end else begin
                  active_thread[(830*4)]   <= 1'b1;
                  active_thread[(830*4)+1] <= 1'b1;
                  active_thread[(830*4)+2] <= 1'b1;
                  active_thread[(830*4)+3] <= 1'b1;
                  spc830_inst_done         <= `ARIANE_CORE830.piton_pc_vld;
                  spc830_phy_pc_w          <= `ARIANE_CORE830.piton_pc;
                end
            end
    

            assign spc831_thread_id = 2'b00;
            assign spc831_rtl_pc = spc831_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(831*4)]   <= 1'b0;
                  active_thread[(831*4)+1] <= 1'b0;
                  active_thread[(831*4)+2] <= 1'b0;
                  active_thread[(831*4)+3] <= 1'b0;
                  spc831_inst_done         <= 0;
                  spc831_phy_pc_w          <= 0;
                end else begin
                  active_thread[(831*4)]   <= 1'b1;
                  active_thread[(831*4)+1] <= 1'b1;
                  active_thread[(831*4)+2] <= 1'b1;
                  active_thread[(831*4)+3] <= 1'b1;
                  spc831_inst_done         <= `ARIANE_CORE831.piton_pc_vld;
                  spc831_phy_pc_w          <= `ARIANE_CORE831.piton_pc;
                end
            end
    

            assign spc832_thread_id = 2'b00;
            assign spc832_rtl_pc = spc832_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(832*4)]   <= 1'b0;
                  active_thread[(832*4)+1] <= 1'b0;
                  active_thread[(832*4)+2] <= 1'b0;
                  active_thread[(832*4)+3] <= 1'b0;
                  spc832_inst_done         <= 0;
                  spc832_phy_pc_w          <= 0;
                end else begin
                  active_thread[(832*4)]   <= 1'b1;
                  active_thread[(832*4)+1] <= 1'b1;
                  active_thread[(832*4)+2] <= 1'b1;
                  active_thread[(832*4)+3] <= 1'b1;
                  spc832_inst_done         <= `ARIANE_CORE832.piton_pc_vld;
                  spc832_phy_pc_w          <= `ARIANE_CORE832.piton_pc;
                end
            end
    

            assign spc833_thread_id = 2'b00;
            assign spc833_rtl_pc = spc833_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(833*4)]   <= 1'b0;
                  active_thread[(833*4)+1] <= 1'b0;
                  active_thread[(833*4)+2] <= 1'b0;
                  active_thread[(833*4)+3] <= 1'b0;
                  spc833_inst_done         <= 0;
                  spc833_phy_pc_w          <= 0;
                end else begin
                  active_thread[(833*4)]   <= 1'b1;
                  active_thread[(833*4)+1] <= 1'b1;
                  active_thread[(833*4)+2] <= 1'b1;
                  active_thread[(833*4)+3] <= 1'b1;
                  spc833_inst_done         <= `ARIANE_CORE833.piton_pc_vld;
                  spc833_phy_pc_w          <= `ARIANE_CORE833.piton_pc;
                end
            end
    

            assign spc834_thread_id = 2'b00;
            assign spc834_rtl_pc = spc834_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(834*4)]   <= 1'b0;
                  active_thread[(834*4)+1] <= 1'b0;
                  active_thread[(834*4)+2] <= 1'b0;
                  active_thread[(834*4)+3] <= 1'b0;
                  spc834_inst_done         <= 0;
                  spc834_phy_pc_w          <= 0;
                end else begin
                  active_thread[(834*4)]   <= 1'b1;
                  active_thread[(834*4)+1] <= 1'b1;
                  active_thread[(834*4)+2] <= 1'b1;
                  active_thread[(834*4)+3] <= 1'b1;
                  spc834_inst_done         <= `ARIANE_CORE834.piton_pc_vld;
                  spc834_phy_pc_w          <= `ARIANE_CORE834.piton_pc;
                end
            end
    

            assign spc835_thread_id = 2'b00;
            assign spc835_rtl_pc = spc835_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(835*4)]   <= 1'b0;
                  active_thread[(835*4)+1] <= 1'b0;
                  active_thread[(835*4)+2] <= 1'b0;
                  active_thread[(835*4)+3] <= 1'b0;
                  spc835_inst_done         <= 0;
                  spc835_phy_pc_w          <= 0;
                end else begin
                  active_thread[(835*4)]   <= 1'b1;
                  active_thread[(835*4)+1] <= 1'b1;
                  active_thread[(835*4)+2] <= 1'b1;
                  active_thread[(835*4)+3] <= 1'b1;
                  spc835_inst_done         <= `ARIANE_CORE835.piton_pc_vld;
                  spc835_phy_pc_w          <= `ARIANE_CORE835.piton_pc;
                end
            end
    

            assign spc836_thread_id = 2'b00;
            assign spc836_rtl_pc = spc836_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(836*4)]   <= 1'b0;
                  active_thread[(836*4)+1] <= 1'b0;
                  active_thread[(836*4)+2] <= 1'b0;
                  active_thread[(836*4)+3] <= 1'b0;
                  spc836_inst_done         <= 0;
                  spc836_phy_pc_w          <= 0;
                end else begin
                  active_thread[(836*4)]   <= 1'b1;
                  active_thread[(836*4)+1] <= 1'b1;
                  active_thread[(836*4)+2] <= 1'b1;
                  active_thread[(836*4)+3] <= 1'b1;
                  spc836_inst_done         <= `ARIANE_CORE836.piton_pc_vld;
                  spc836_phy_pc_w          <= `ARIANE_CORE836.piton_pc;
                end
            end
    

            assign spc837_thread_id = 2'b00;
            assign spc837_rtl_pc = spc837_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(837*4)]   <= 1'b0;
                  active_thread[(837*4)+1] <= 1'b0;
                  active_thread[(837*4)+2] <= 1'b0;
                  active_thread[(837*4)+3] <= 1'b0;
                  spc837_inst_done         <= 0;
                  spc837_phy_pc_w          <= 0;
                end else begin
                  active_thread[(837*4)]   <= 1'b1;
                  active_thread[(837*4)+1] <= 1'b1;
                  active_thread[(837*4)+2] <= 1'b1;
                  active_thread[(837*4)+3] <= 1'b1;
                  spc837_inst_done         <= `ARIANE_CORE837.piton_pc_vld;
                  spc837_phy_pc_w          <= `ARIANE_CORE837.piton_pc;
                end
            end
    

            assign spc838_thread_id = 2'b00;
            assign spc838_rtl_pc = spc838_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(838*4)]   <= 1'b0;
                  active_thread[(838*4)+1] <= 1'b0;
                  active_thread[(838*4)+2] <= 1'b0;
                  active_thread[(838*4)+3] <= 1'b0;
                  spc838_inst_done         <= 0;
                  spc838_phy_pc_w          <= 0;
                end else begin
                  active_thread[(838*4)]   <= 1'b1;
                  active_thread[(838*4)+1] <= 1'b1;
                  active_thread[(838*4)+2] <= 1'b1;
                  active_thread[(838*4)+3] <= 1'b1;
                  spc838_inst_done         <= `ARIANE_CORE838.piton_pc_vld;
                  spc838_phy_pc_w          <= `ARIANE_CORE838.piton_pc;
                end
            end
    

            assign spc839_thread_id = 2'b00;
            assign spc839_rtl_pc = spc839_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(839*4)]   <= 1'b0;
                  active_thread[(839*4)+1] <= 1'b0;
                  active_thread[(839*4)+2] <= 1'b0;
                  active_thread[(839*4)+3] <= 1'b0;
                  spc839_inst_done         <= 0;
                  spc839_phy_pc_w          <= 0;
                end else begin
                  active_thread[(839*4)]   <= 1'b1;
                  active_thread[(839*4)+1] <= 1'b1;
                  active_thread[(839*4)+2] <= 1'b1;
                  active_thread[(839*4)+3] <= 1'b1;
                  spc839_inst_done         <= `ARIANE_CORE839.piton_pc_vld;
                  spc839_phy_pc_w          <= `ARIANE_CORE839.piton_pc;
                end
            end
    

            assign spc840_thread_id = 2'b00;
            assign spc840_rtl_pc = spc840_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(840*4)]   <= 1'b0;
                  active_thread[(840*4)+1] <= 1'b0;
                  active_thread[(840*4)+2] <= 1'b0;
                  active_thread[(840*4)+3] <= 1'b0;
                  spc840_inst_done         <= 0;
                  spc840_phy_pc_w          <= 0;
                end else begin
                  active_thread[(840*4)]   <= 1'b1;
                  active_thread[(840*4)+1] <= 1'b1;
                  active_thread[(840*4)+2] <= 1'b1;
                  active_thread[(840*4)+3] <= 1'b1;
                  spc840_inst_done         <= `ARIANE_CORE840.piton_pc_vld;
                  spc840_phy_pc_w          <= `ARIANE_CORE840.piton_pc;
                end
            end
    

            assign spc841_thread_id = 2'b00;
            assign spc841_rtl_pc = spc841_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(841*4)]   <= 1'b0;
                  active_thread[(841*4)+1] <= 1'b0;
                  active_thread[(841*4)+2] <= 1'b0;
                  active_thread[(841*4)+3] <= 1'b0;
                  spc841_inst_done         <= 0;
                  spc841_phy_pc_w          <= 0;
                end else begin
                  active_thread[(841*4)]   <= 1'b1;
                  active_thread[(841*4)+1] <= 1'b1;
                  active_thread[(841*4)+2] <= 1'b1;
                  active_thread[(841*4)+3] <= 1'b1;
                  spc841_inst_done         <= `ARIANE_CORE841.piton_pc_vld;
                  spc841_phy_pc_w          <= `ARIANE_CORE841.piton_pc;
                end
            end
    

            assign spc842_thread_id = 2'b00;
            assign spc842_rtl_pc = spc842_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(842*4)]   <= 1'b0;
                  active_thread[(842*4)+1] <= 1'b0;
                  active_thread[(842*4)+2] <= 1'b0;
                  active_thread[(842*4)+3] <= 1'b0;
                  spc842_inst_done         <= 0;
                  spc842_phy_pc_w          <= 0;
                end else begin
                  active_thread[(842*4)]   <= 1'b1;
                  active_thread[(842*4)+1] <= 1'b1;
                  active_thread[(842*4)+2] <= 1'b1;
                  active_thread[(842*4)+3] <= 1'b1;
                  spc842_inst_done         <= `ARIANE_CORE842.piton_pc_vld;
                  spc842_phy_pc_w          <= `ARIANE_CORE842.piton_pc;
                end
            end
    

            assign spc843_thread_id = 2'b00;
            assign spc843_rtl_pc = spc843_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(843*4)]   <= 1'b0;
                  active_thread[(843*4)+1] <= 1'b0;
                  active_thread[(843*4)+2] <= 1'b0;
                  active_thread[(843*4)+3] <= 1'b0;
                  spc843_inst_done         <= 0;
                  spc843_phy_pc_w          <= 0;
                end else begin
                  active_thread[(843*4)]   <= 1'b1;
                  active_thread[(843*4)+1] <= 1'b1;
                  active_thread[(843*4)+2] <= 1'b1;
                  active_thread[(843*4)+3] <= 1'b1;
                  spc843_inst_done         <= `ARIANE_CORE843.piton_pc_vld;
                  spc843_phy_pc_w          <= `ARIANE_CORE843.piton_pc;
                end
            end
    

            assign spc844_thread_id = 2'b00;
            assign spc844_rtl_pc = spc844_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(844*4)]   <= 1'b0;
                  active_thread[(844*4)+1] <= 1'b0;
                  active_thread[(844*4)+2] <= 1'b0;
                  active_thread[(844*4)+3] <= 1'b0;
                  spc844_inst_done         <= 0;
                  spc844_phy_pc_w          <= 0;
                end else begin
                  active_thread[(844*4)]   <= 1'b1;
                  active_thread[(844*4)+1] <= 1'b1;
                  active_thread[(844*4)+2] <= 1'b1;
                  active_thread[(844*4)+3] <= 1'b1;
                  spc844_inst_done         <= `ARIANE_CORE844.piton_pc_vld;
                  spc844_phy_pc_w          <= `ARIANE_CORE844.piton_pc;
                end
            end
    

            assign spc845_thread_id = 2'b00;
            assign spc845_rtl_pc = spc845_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(845*4)]   <= 1'b0;
                  active_thread[(845*4)+1] <= 1'b0;
                  active_thread[(845*4)+2] <= 1'b0;
                  active_thread[(845*4)+3] <= 1'b0;
                  spc845_inst_done         <= 0;
                  spc845_phy_pc_w          <= 0;
                end else begin
                  active_thread[(845*4)]   <= 1'b1;
                  active_thread[(845*4)+1] <= 1'b1;
                  active_thread[(845*4)+2] <= 1'b1;
                  active_thread[(845*4)+3] <= 1'b1;
                  spc845_inst_done         <= `ARIANE_CORE845.piton_pc_vld;
                  spc845_phy_pc_w          <= `ARIANE_CORE845.piton_pc;
                end
            end
    

            assign spc846_thread_id = 2'b00;
            assign spc846_rtl_pc = spc846_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(846*4)]   <= 1'b0;
                  active_thread[(846*4)+1] <= 1'b0;
                  active_thread[(846*4)+2] <= 1'b0;
                  active_thread[(846*4)+3] <= 1'b0;
                  spc846_inst_done         <= 0;
                  spc846_phy_pc_w          <= 0;
                end else begin
                  active_thread[(846*4)]   <= 1'b1;
                  active_thread[(846*4)+1] <= 1'b1;
                  active_thread[(846*4)+2] <= 1'b1;
                  active_thread[(846*4)+3] <= 1'b1;
                  spc846_inst_done         <= `ARIANE_CORE846.piton_pc_vld;
                  spc846_phy_pc_w          <= `ARIANE_CORE846.piton_pc;
                end
            end
    

            assign spc847_thread_id = 2'b00;
            assign spc847_rtl_pc = spc847_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(847*4)]   <= 1'b0;
                  active_thread[(847*4)+1] <= 1'b0;
                  active_thread[(847*4)+2] <= 1'b0;
                  active_thread[(847*4)+3] <= 1'b0;
                  spc847_inst_done         <= 0;
                  spc847_phy_pc_w          <= 0;
                end else begin
                  active_thread[(847*4)]   <= 1'b1;
                  active_thread[(847*4)+1] <= 1'b1;
                  active_thread[(847*4)+2] <= 1'b1;
                  active_thread[(847*4)+3] <= 1'b1;
                  spc847_inst_done         <= `ARIANE_CORE847.piton_pc_vld;
                  spc847_phy_pc_w          <= `ARIANE_CORE847.piton_pc;
                end
            end
    

            assign spc848_thread_id = 2'b00;
            assign spc848_rtl_pc = spc848_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(848*4)]   <= 1'b0;
                  active_thread[(848*4)+1] <= 1'b0;
                  active_thread[(848*4)+2] <= 1'b0;
                  active_thread[(848*4)+3] <= 1'b0;
                  spc848_inst_done         <= 0;
                  spc848_phy_pc_w          <= 0;
                end else begin
                  active_thread[(848*4)]   <= 1'b1;
                  active_thread[(848*4)+1] <= 1'b1;
                  active_thread[(848*4)+2] <= 1'b1;
                  active_thread[(848*4)+3] <= 1'b1;
                  spc848_inst_done         <= `ARIANE_CORE848.piton_pc_vld;
                  spc848_phy_pc_w          <= `ARIANE_CORE848.piton_pc;
                end
            end
    

            assign spc849_thread_id = 2'b00;
            assign spc849_rtl_pc = spc849_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(849*4)]   <= 1'b0;
                  active_thread[(849*4)+1] <= 1'b0;
                  active_thread[(849*4)+2] <= 1'b0;
                  active_thread[(849*4)+3] <= 1'b0;
                  spc849_inst_done         <= 0;
                  spc849_phy_pc_w          <= 0;
                end else begin
                  active_thread[(849*4)]   <= 1'b1;
                  active_thread[(849*4)+1] <= 1'b1;
                  active_thread[(849*4)+2] <= 1'b1;
                  active_thread[(849*4)+3] <= 1'b1;
                  spc849_inst_done         <= `ARIANE_CORE849.piton_pc_vld;
                  spc849_phy_pc_w          <= `ARIANE_CORE849.piton_pc;
                end
            end
    

            assign spc850_thread_id = 2'b00;
            assign spc850_rtl_pc = spc850_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(850*4)]   <= 1'b0;
                  active_thread[(850*4)+1] <= 1'b0;
                  active_thread[(850*4)+2] <= 1'b0;
                  active_thread[(850*4)+3] <= 1'b0;
                  spc850_inst_done         <= 0;
                  spc850_phy_pc_w          <= 0;
                end else begin
                  active_thread[(850*4)]   <= 1'b1;
                  active_thread[(850*4)+1] <= 1'b1;
                  active_thread[(850*4)+2] <= 1'b1;
                  active_thread[(850*4)+3] <= 1'b1;
                  spc850_inst_done         <= `ARIANE_CORE850.piton_pc_vld;
                  spc850_phy_pc_w          <= `ARIANE_CORE850.piton_pc;
                end
            end
    

            assign spc851_thread_id = 2'b00;
            assign spc851_rtl_pc = spc851_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(851*4)]   <= 1'b0;
                  active_thread[(851*4)+1] <= 1'b0;
                  active_thread[(851*4)+2] <= 1'b0;
                  active_thread[(851*4)+3] <= 1'b0;
                  spc851_inst_done         <= 0;
                  spc851_phy_pc_w          <= 0;
                end else begin
                  active_thread[(851*4)]   <= 1'b1;
                  active_thread[(851*4)+1] <= 1'b1;
                  active_thread[(851*4)+2] <= 1'b1;
                  active_thread[(851*4)+3] <= 1'b1;
                  spc851_inst_done         <= `ARIANE_CORE851.piton_pc_vld;
                  spc851_phy_pc_w          <= `ARIANE_CORE851.piton_pc;
                end
            end
    

            assign spc852_thread_id = 2'b00;
            assign spc852_rtl_pc = spc852_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(852*4)]   <= 1'b0;
                  active_thread[(852*4)+1] <= 1'b0;
                  active_thread[(852*4)+2] <= 1'b0;
                  active_thread[(852*4)+3] <= 1'b0;
                  spc852_inst_done         <= 0;
                  spc852_phy_pc_w          <= 0;
                end else begin
                  active_thread[(852*4)]   <= 1'b1;
                  active_thread[(852*4)+1] <= 1'b1;
                  active_thread[(852*4)+2] <= 1'b1;
                  active_thread[(852*4)+3] <= 1'b1;
                  spc852_inst_done         <= `ARIANE_CORE852.piton_pc_vld;
                  spc852_phy_pc_w          <= `ARIANE_CORE852.piton_pc;
                end
            end
    

            assign spc853_thread_id = 2'b00;
            assign spc853_rtl_pc = spc853_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(853*4)]   <= 1'b0;
                  active_thread[(853*4)+1] <= 1'b0;
                  active_thread[(853*4)+2] <= 1'b0;
                  active_thread[(853*4)+3] <= 1'b0;
                  spc853_inst_done         <= 0;
                  spc853_phy_pc_w          <= 0;
                end else begin
                  active_thread[(853*4)]   <= 1'b1;
                  active_thread[(853*4)+1] <= 1'b1;
                  active_thread[(853*4)+2] <= 1'b1;
                  active_thread[(853*4)+3] <= 1'b1;
                  spc853_inst_done         <= `ARIANE_CORE853.piton_pc_vld;
                  spc853_phy_pc_w          <= `ARIANE_CORE853.piton_pc;
                end
            end
    

            assign spc854_thread_id = 2'b00;
            assign spc854_rtl_pc = spc854_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(854*4)]   <= 1'b0;
                  active_thread[(854*4)+1] <= 1'b0;
                  active_thread[(854*4)+2] <= 1'b0;
                  active_thread[(854*4)+3] <= 1'b0;
                  spc854_inst_done         <= 0;
                  spc854_phy_pc_w          <= 0;
                end else begin
                  active_thread[(854*4)]   <= 1'b1;
                  active_thread[(854*4)+1] <= 1'b1;
                  active_thread[(854*4)+2] <= 1'b1;
                  active_thread[(854*4)+3] <= 1'b1;
                  spc854_inst_done         <= `ARIANE_CORE854.piton_pc_vld;
                  spc854_phy_pc_w          <= `ARIANE_CORE854.piton_pc;
                end
            end
    

            assign spc855_thread_id = 2'b00;
            assign spc855_rtl_pc = spc855_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(855*4)]   <= 1'b0;
                  active_thread[(855*4)+1] <= 1'b0;
                  active_thread[(855*4)+2] <= 1'b0;
                  active_thread[(855*4)+3] <= 1'b0;
                  spc855_inst_done         <= 0;
                  spc855_phy_pc_w          <= 0;
                end else begin
                  active_thread[(855*4)]   <= 1'b1;
                  active_thread[(855*4)+1] <= 1'b1;
                  active_thread[(855*4)+2] <= 1'b1;
                  active_thread[(855*4)+3] <= 1'b1;
                  spc855_inst_done         <= `ARIANE_CORE855.piton_pc_vld;
                  spc855_phy_pc_w          <= `ARIANE_CORE855.piton_pc;
                end
            end
    

            assign spc856_thread_id = 2'b00;
            assign spc856_rtl_pc = spc856_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(856*4)]   <= 1'b0;
                  active_thread[(856*4)+1] <= 1'b0;
                  active_thread[(856*4)+2] <= 1'b0;
                  active_thread[(856*4)+3] <= 1'b0;
                  spc856_inst_done         <= 0;
                  spc856_phy_pc_w          <= 0;
                end else begin
                  active_thread[(856*4)]   <= 1'b1;
                  active_thread[(856*4)+1] <= 1'b1;
                  active_thread[(856*4)+2] <= 1'b1;
                  active_thread[(856*4)+3] <= 1'b1;
                  spc856_inst_done         <= `ARIANE_CORE856.piton_pc_vld;
                  spc856_phy_pc_w          <= `ARIANE_CORE856.piton_pc;
                end
            end
    

            assign spc857_thread_id = 2'b00;
            assign spc857_rtl_pc = spc857_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(857*4)]   <= 1'b0;
                  active_thread[(857*4)+1] <= 1'b0;
                  active_thread[(857*4)+2] <= 1'b0;
                  active_thread[(857*4)+3] <= 1'b0;
                  spc857_inst_done         <= 0;
                  spc857_phy_pc_w          <= 0;
                end else begin
                  active_thread[(857*4)]   <= 1'b1;
                  active_thread[(857*4)+1] <= 1'b1;
                  active_thread[(857*4)+2] <= 1'b1;
                  active_thread[(857*4)+3] <= 1'b1;
                  spc857_inst_done         <= `ARIANE_CORE857.piton_pc_vld;
                  spc857_phy_pc_w          <= `ARIANE_CORE857.piton_pc;
                end
            end
    

            assign spc858_thread_id = 2'b00;
            assign spc858_rtl_pc = spc858_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(858*4)]   <= 1'b0;
                  active_thread[(858*4)+1] <= 1'b0;
                  active_thread[(858*4)+2] <= 1'b0;
                  active_thread[(858*4)+3] <= 1'b0;
                  spc858_inst_done         <= 0;
                  spc858_phy_pc_w          <= 0;
                end else begin
                  active_thread[(858*4)]   <= 1'b1;
                  active_thread[(858*4)+1] <= 1'b1;
                  active_thread[(858*4)+2] <= 1'b1;
                  active_thread[(858*4)+3] <= 1'b1;
                  spc858_inst_done         <= `ARIANE_CORE858.piton_pc_vld;
                  spc858_phy_pc_w          <= `ARIANE_CORE858.piton_pc;
                end
            end
    

            assign spc859_thread_id = 2'b00;
            assign spc859_rtl_pc = spc859_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(859*4)]   <= 1'b0;
                  active_thread[(859*4)+1] <= 1'b0;
                  active_thread[(859*4)+2] <= 1'b0;
                  active_thread[(859*4)+3] <= 1'b0;
                  spc859_inst_done         <= 0;
                  spc859_phy_pc_w          <= 0;
                end else begin
                  active_thread[(859*4)]   <= 1'b1;
                  active_thread[(859*4)+1] <= 1'b1;
                  active_thread[(859*4)+2] <= 1'b1;
                  active_thread[(859*4)+3] <= 1'b1;
                  spc859_inst_done         <= `ARIANE_CORE859.piton_pc_vld;
                  spc859_phy_pc_w          <= `ARIANE_CORE859.piton_pc;
                end
            end
    

            assign spc860_thread_id = 2'b00;
            assign spc860_rtl_pc = spc860_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(860*4)]   <= 1'b0;
                  active_thread[(860*4)+1] <= 1'b0;
                  active_thread[(860*4)+2] <= 1'b0;
                  active_thread[(860*4)+3] <= 1'b0;
                  spc860_inst_done         <= 0;
                  spc860_phy_pc_w          <= 0;
                end else begin
                  active_thread[(860*4)]   <= 1'b1;
                  active_thread[(860*4)+1] <= 1'b1;
                  active_thread[(860*4)+2] <= 1'b1;
                  active_thread[(860*4)+3] <= 1'b1;
                  spc860_inst_done         <= `ARIANE_CORE860.piton_pc_vld;
                  spc860_phy_pc_w          <= `ARIANE_CORE860.piton_pc;
                end
            end
    

            assign spc861_thread_id = 2'b00;
            assign spc861_rtl_pc = spc861_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(861*4)]   <= 1'b0;
                  active_thread[(861*4)+1] <= 1'b0;
                  active_thread[(861*4)+2] <= 1'b0;
                  active_thread[(861*4)+3] <= 1'b0;
                  spc861_inst_done         <= 0;
                  spc861_phy_pc_w          <= 0;
                end else begin
                  active_thread[(861*4)]   <= 1'b1;
                  active_thread[(861*4)+1] <= 1'b1;
                  active_thread[(861*4)+2] <= 1'b1;
                  active_thread[(861*4)+3] <= 1'b1;
                  spc861_inst_done         <= `ARIANE_CORE861.piton_pc_vld;
                  spc861_phy_pc_w          <= `ARIANE_CORE861.piton_pc;
                end
            end
    

            assign spc862_thread_id = 2'b00;
            assign spc862_rtl_pc = spc862_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(862*4)]   <= 1'b0;
                  active_thread[(862*4)+1] <= 1'b0;
                  active_thread[(862*4)+2] <= 1'b0;
                  active_thread[(862*4)+3] <= 1'b0;
                  spc862_inst_done         <= 0;
                  spc862_phy_pc_w          <= 0;
                end else begin
                  active_thread[(862*4)]   <= 1'b1;
                  active_thread[(862*4)+1] <= 1'b1;
                  active_thread[(862*4)+2] <= 1'b1;
                  active_thread[(862*4)+3] <= 1'b1;
                  spc862_inst_done         <= `ARIANE_CORE862.piton_pc_vld;
                  spc862_phy_pc_w          <= `ARIANE_CORE862.piton_pc;
                end
            end
    

            assign spc863_thread_id = 2'b00;
            assign spc863_rtl_pc = spc863_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(863*4)]   <= 1'b0;
                  active_thread[(863*4)+1] <= 1'b0;
                  active_thread[(863*4)+2] <= 1'b0;
                  active_thread[(863*4)+3] <= 1'b0;
                  spc863_inst_done         <= 0;
                  spc863_phy_pc_w          <= 0;
                end else begin
                  active_thread[(863*4)]   <= 1'b1;
                  active_thread[(863*4)+1] <= 1'b1;
                  active_thread[(863*4)+2] <= 1'b1;
                  active_thread[(863*4)+3] <= 1'b1;
                  spc863_inst_done         <= `ARIANE_CORE863.piton_pc_vld;
                  spc863_phy_pc_w          <= `ARIANE_CORE863.piton_pc;
                end
            end
    

            assign spc864_thread_id = 2'b00;
            assign spc864_rtl_pc = spc864_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(864*4)]   <= 1'b0;
                  active_thread[(864*4)+1] <= 1'b0;
                  active_thread[(864*4)+2] <= 1'b0;
                  active_thread[(864*4)+3] <= 1'b0;
                  spc864_inst_done         <= 0;
                  spc864_phy_pc_w          <= 0;
                end else begin
                  active_thread[(864*4)]   <= 1'b1;
                  active_thread[(864*4)+1] <= 1'b1;
                  active_thread[(864*4)+2] <= 1'b1;
                  active_thread[(864*4)+3] <= 1'b1;
                  spc864_inst_done         <= `ARIANE_CORE864.piton_pc_vld;
                  spc864_phy_pc_w          <= `ARIANE_CORE864.piton_pc;
                end
            end
    

            assign spc865_thread_id = 2'b00;
            assign spc865_rtl_pc = spc865_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(865*4)]   <= 1'b0;
                  active_thread[(865*4)+1] <= 1'b0;
                  active_thread[(865*4)+2] <= 1'b0;
                  active_thread[(865*4)+3] <= 1'b0;
                  spc865_inst_done         <= 0;
                  spc865_phy_pc_w          <= 0;
                end else begin
                  active_thread[(865*4)]   <= 1'b1;
                  active_thread[(865*4)+1] <= 1'b1;
                  active_thread[(865*4)+2] <= 1'b1;
                  active_thread[(865*4)+3] <= 1'b1;
                  spc865_inst_done         <= `ARIANE_CORE865.piton_pc_vld;
                  spc865_phy_pc_w          <= `ARIANE_CORE865.piton_pc;
                end
            end
    

            assign spc866_thread_id = 2'b00;
            assign spc866_rtl_pc = spc866_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(866*4)]   <= 1'b0;
                  active_thread[(866*4)+1] <= 1'b0;
                  active_thread[(866*4)+2] <= 1'b0;
                  active_thread[(866*4)+3] <= 1'b0;
                  spc866_inst_done         <= 0;
                  spc866_phy_pc_w          <= 0;
                end else begin
                  active_thread[(866*4)]   <= 1'b1;
                  active_thread[(866*4)+1] <= 1'b1;
                  active_thread[(866*4)+2] <= 1'b1;
                  active_thread[(866*4)+3] <= 1'b1;
                  spc866_inst_done         <= `ARIANE_CORE866.piton_pc_vld;
                  spc866_phy_pc_w          <= `ARIANE_CORE866.piton_pc;
                end
            end
    

            assign spc867_thread_id = 2'b00;
            assign spc867_rtl_pc = spc867_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(867*4)]   <= 1'b0;
                  active_thread[(867*4)+1] <= 1'b0;
                  active_thread[(867*4)+2] <= 1'b0;
                  active_thread[(867*4)+3] <= 1'b0;
                  spc867_inst_done         <= 0;
                  spc867_phy_pc_w          <= 0;
                end else begin
                  active_thread[(867*4)]   <= 1'b1;
                  active_thread[(867*4)+1] <= 1'b1;
                  active_thread[(867*4)+2] <= 1'b1;
                  active_thread[(867*4)+3] <= 1'b1;
                  spc867_inst_done         <= `ARIANE_CORE867.piton_pc_vld;
                  spc867_phy_pc_w          <= `ARIANE_CORE867.piton_pc;
                end
            end
    

            assign spc868_thread_id = 2'b00;
            assign spc868_rtl_pc = spc868_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(868*4)]   <= 1'b0;
                  active_thread[(868*4)+1] <= 1'b0;
                  active_thread[(868*4)+2] <= 1'b0;
                  active_thread[(868*4)+3] <= 1'b0;
                  spc868_inst_done         <= 0;
                  spc868_phy_pc_w          <= 0;
                end else begin
                  active_thread[(868*4)]   <= 1'b1;
                  active_thread[(868*4)+1] <= 1'b1;
                  active_thread[(868*4)+2] <= 1'b1;
                  active_thread[(868*4)+3] <= 1'b1;
                  spc868_inst_done         <= `ARIANE_CORE868.piton_pc_vld;
                  spc868_phy_pc_w          <= `ARIANE_CORE868.piton_pc;
                end
            end
    

            assign spc869_thread_id = 2'b00;
            assign spc869_rtl_pc = spc869_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(869*4)]   <= 1'b0;
                  active_thread[(869*4)+1] <= 1'b0;
                  active_thread[(869*4)+2] <= 1'b0;
                  active_thread[(869*4)+3] <= 1'b0;
                  spc869_inst_done         <= 0;
                  spc869_phy_pc_w          <= 0;
                end else begin
                  active_thread[(869*4)]   <= 1'b1;
                  active_thread[(869*4)+1] <= 1'b1;
                  active_thread[(869*4)+2] <= 1'b1;
                  active_thread[(869*4)+3] <= 1'b1;
                  spc869_inst_done         <= `ARIANE_CORE869.piton_pc_vld;
                  spc869_phy_pc_w          <= `ARIANE_CORE869.piton_pc;
                end
            end
    

            assign spc870_thread_id = 2'b00;
            assign spc870_rtl_pc = spc870_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(870*4)]   <= 1'b0;
                  active_thread[(870*4)+1] <= 1'b0;
                  active_thread[(870*4)+2] <= 1'b0;
                  active_thread[(870*4)+3] <= 1'b0;
                  spc870_inst_done         <= 0;
                  spc870_phy_pc_w          <= 0;
                end else begin
                  active_thread[(870*4)]   <= 1'b1;
                  active_thread[(870*4)+1] <= 1'b1;
                  active_thread[(870*4)+2] <= 1'b1;
                  active_thread[(870*4)+3] <= 1'b1;
                  spc870_inst_done         <= `ARIANE_CORE870.piton_pc_vld;
                  spc870_phy_pc_w          <= `ARIANE_CORE870.piton_pc;
                end
            end
    

            assign spc871_thread_id = 2'b00;
            assign spc871_rtl_pc = spc871_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(871*4)]   <= 1'b0;
                  active_thread[(871*4)+1] <= 1'b0;
                  active_thread[(871*4)+2] <= 1'b0;
                  active_thread[(871*4)+3] <= 1'b0;
                  spc871_inst_done         <= 0;
                  spc871_phy_pc_w          <= 0;
                end else begin
                  active_thread[(871*4)]   <= 1'b1;
                  active_thread[(871*4)+1] <= 1'b1;
                  active_thread[(871*4)+2] <= 1'b1;
                  active_thread[(871*4)+3] <= 1'b1;
                  spc871_inst_done         <= `ARIANE_CORE871.piton_pc_vld;
                  spc871_phy_pc_w          <= `ARIANE_CORE871.piton_pc;
                end
            end
    

            assign spc872_thread_id = 2'b00;
            assign spc872_rtl_pc = spc872_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(872*4)]   <= 1'b0;
                  active_thread[(872*4)+1] <= 1'b0;
                  active_thread[(872*4)+2] <= 1'b0;
                  active_thread[(872*4)+3] <= 1'b0;
                  spc872_inst_done         <= 0;
                  spc872_phy_pc_w          <= 0;
                end else begin
                  active_thread[(872*4)]   <= 1'b1;
                  active_thread[(872*4)+1] <= 1'b1;
                  active_thread[(872*4)+2] <= 1'b1;
                  active_thread[(872*4)+3] <= 1'b1;
                  spc872_inst_done         <= `ARIANE_CORE872.piton_pc_vld;
                  spc872_phy_pc_w          <= `ARIANE_CORE872.piton_pc;
                end
            end
    

            assign spc873_thread_id = 2'b00;
            assign spc873_rtl_pc = spc873_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(873*4)]   <= 1'b0;
                  active_thread[(873*4)+1] <= 1'b0;
                  active_thread[(873*4)+2] <= 1'b0;
                  active_thread[(873*4)+3] <= 1'b0;
                  spc873_inst_done         <= 0;
                  spc873_phy_pc_w          <= 0;
                end else begin
                  active_thread[(873*4)]   <= 1'b1;
                  active_thread[(873*4)+1] <= 1'b1;
                  active_thread[(873*4)+2] <= 1'b1;
                  active_thread[(873*4)+3] <= 1'b1;
                  spc873_inst_done         <= `ARIANE_CORE873.piton_pc_vld;
                  spc873_phy_pc_w          <= `ARIANE_CORE873.piton_pc;
                end
            end
    

            assign spc874_thread_id = 2'b00;
            assign spc874_rtl_pc = spc874_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(874*4)]   <= 1'b0;
                  active_thread[(874*4)+1] <= 1'b0;
                  active_thread[(874*4)+2] <= 1'b0;
                  active_thread[(874*4)+3] <= 1'b0;
                  spc874_inst_done         <= 0;
                  spc874_phy_pc_w          <= 0;
                end else begin
                  active_thread[(874*4)]   <= 1'b1;
                  active_thread[(874*4)+1] <= 1'b1;
                  active_thread[(874*4)+2] <= 1'b1;
                  active_thread[(874*4)+3] <= 1'b1;
                  spc874_inst_done         <= `ARIANE_CORE874.piton_pc_vld;
                  spc874_phy_pc_w          <= `ARIANE_CORE874.piton_pc;
                end
            end
    

            assign spc875_thread_id = 2'b00;
            assign spc875_rtl_pc = spc875_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(875*4)]   <= 1'b0;
                  active_thread[(875*4)+1] <= 1'b0;
                  active_thread[(875*4)+2] <= 1'b0;
                  active_thread[(875*4)+3] <= 1'b0;
                  spc875_inst_done         <= 0;
                  spc875_phy_pc_w          <= 0;
                end else begin
                  active_thread[(875*4)]   <= 1'b1;
                  active_thread[(875*4)+1] <= 1'b1;
                  active_thread[(875*4)+2] <= 1'b1;
                  active_thread[(875*4)+3] <= 1'b1;
                  spc875_inst_done         <= `ARIANE_CORE875.piton_pc_vld;
                  spc875_phy_pc_w          <= `ARIANE_CORE875.piton_pc;
                end
            end
    

            assign spc876_thread_id = 2'b00;
            assign spc876_rtl_pc = spc876_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(876*4)]   <= 1'b0;
                  active_thread[(876*4)+1] <= 1'b0;
                  active_thread[(876*4)+2] <= 1'b0;
                  active_thread[(876*4)+3] <= 1'b0;
                  spc876_inst_done         <= 0;
                  spc876_phy_pc_w          <= 0;
                end else begin
                  active_thread[(876*4)]   <= 1'b1;
                  active_thread[(876*4)+1] <= 1'b1;
                  active_thread[(876*4)+2] <= 1'b1;
                  active_thread[(876*4)+3] <= 1'b1;
                  spc876_inst_done         <= `ARIANE_CORE876.piton_pc_vld;
                  spc876_phy_pc_w          <= `ARIANE_CORE876.piton_pc;
                end
            end
    

            assign spc877_thread_id = 2'b00;
            assign spc877_rtl_pc = spc877_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(877*4)]   <= 1'b0;
                  active_thread[(877*4)+1] <= 1'b0;
                  active_thread[(877*4)+2] <= 1'b0;
                  active_thread[(877*4)+3] <= 1'b0;
                  spc877_inst_done         <= 0;
                  spc877_phy_pc_w          <= 0;
                end else begin
                  active_thread[(877*4)]   <= 1'b1;
                  active_thread[(877*4)+1] <= 1'b1;
                  active_thread[(877*4)+2] <= 1'b1;
                  active_thread[(877*4)+3] <= 1'b1;
                  spc877_inst_done         <= `ARIANE_CORE877.piton_pc_vld;
                  spc877_phy_pc_w          <= `ARIANE_CORE877.piton_pc;
                end
            end
    

            assign spc878_thread_id = 2'b00;
            assign spc878_rtl_pc = spc878_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(878*4)]   <= 1'b0;
                  active_thread[(878*4)+1] <= 1'b0;
                  active_thread[(878*4)+2] <= 1'b0;
                  active_thread[(878*4)+3] <= 1'b0;
                  spc878_inst_done         <= 0;
                  spc878_phy_pc_w          <= 0;
                end else begin
                  active_thread[(878*4)]   <= 1'b1;
                  active_thread[(878*4)+1] <= 1'b1;
                  active_thread[(878*4)+2] <= 1'b1;
                  active_thread[(878*4)+3] <= 1'b1;
                  spc878_inst_done         <= `ARIANE_CORE878.piton_pc_vld;
                  spc878_phy_pc_w          <= `ARIANE_CORE878.piton_pc;
                end
            end
    

            assign spc879_thread_id = 2'b00;
            assign spc879_rtl_pc = spc879_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(879*4)]   <= 1'b0;
                  active_thread[(879*4)+1] <= 1'b0;
                  active_thread[(879*4)+2] <= 1'b0;
                  active_thread[(879*4)+3] <= 1'b0;
                  spc879_inst_done         <= 0;
                  spc879_phy_pc_w          <= 0;
                end else begin
                  active_thread[(879*4)]   <= 1'b1;
                  active_thread[(879*4)+1] <= 1'b1;
                  active_thread[(879*4)+2] <= 1'b1;
                  active_thread[(879*4)+3] <= 1'b1;
                  spc879_inst_done         <= `ARIANE_CORE879.piton_pc_vld;
                  spc879_phy_pc_w          <= `ARIANE_CORE879.piton_pc;
                end
            end
    

            assign spc880_thread_id = 2'b00;
            assign spc880_rtl_pc = spc880_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(880*4)]   <= 1'b0;
                  active_thread[(880*4)+1] <= 1'b0;
                  active_thread[(880*4)+2] <= 1'b0;
                  active_thread[(880*4)+3] <= 1'b0;
                  spc880_inst_done         <= 0;
                  spc880_phy_pc_w          <= 0;
                end else begin
                  active_thread[(880*4)]   <= 1'b1;
                  active_thread[(880*4)+1] <= 1'b1;
                  active_thread[(880*4)+2] <= 1'b1;
                  active_thread[(880*4)+3] <= 1'b1;
                  spc880_inst_done         <= `ARIANE_CORE880.piton_pc_vld;
                  spc880_phy_pc_w          <= `ARIANE_CORE880.piton_pc;
                end
            end
    

            assign spc881_thread_id = 2'b00;
            assign spc881_rtl_pc = spc881_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(881*4)]   <= 1'b0;
                  active_thread[(881*4)+1] <= 1'b0;
                  active_thread[(881*4)+2] <= 1'b0;
                  active_thread[(881*4)+3] <= 1'b0;
                  spc881_inst_done         <= 0;
                  spc881_phy_pc_w          <= 0;
                end else begin
                  active_thread[(881*4)]   <= 1'b1;
                  active_thread[(881*4)+1] <= 1'b1;
                  active_thread[(881*4)+2] <= 1'b1;
                  active_thread[(881*4)+3] <= 1'b1;
                  spc881_inst_done         <= `ARIANE_CORE881.piton_pc_vld;
                  spc881_phy_pc_w          <= `ARIANE_CORE881.piton_pc;
                end
            end
    

            assign spc882_thread_id = 2'b00;
            assign spc882_rtl_pc = spc882_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(882*4)]   <= 1'b0;
                  active_thread[(882*4)+1] <= 1'b0;
                  active_thread[(882*4)+2] <= 1'b0;
                  active_thread[(882*4)+3] <= 1'b0;
                  spc882_inst_done         <= 0;
                  spc882_phy_pc_w          <= 0;
                end else begin
                  active_thread[(882*4)]   <= 1'b1;
                  active_thread[(882*4)+1] <= 1'b1;
                  active_thread[(882*4)+2] <= 1'b1;
                  active_thread[(882*4)+3] <= 1'b1;
                  spc882_inst_done         <= `ARIANE_CORE882.piton_pc_vld;
                  spc882_phy_pc_w          <= `ARIANE_CORE882.piton_pc;
                end
            end
    

            assign spc883_thread_id = 2'b00;
            assign spc883_rtl_pc = spc883_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(883*4)]   <= 1'b0;
                  active_thread[(883*4)+1] <= 1'b0;
                  active_thread[(883*4)+2] <= 1'b0;
                  active_thread[(883*4)+3] <= 1'b0;
                  spc883_inst_done         <= 0;
                  spc883_phy_pc_w          <= 0;
                end else begin
                  active_thread[(883*4)]   <= 1'b1;
                  active_thread[(883*4)+1] <= 1'b1;
                  active_thread[(883*4)+2] <= 1'b1;
                  active_thread[(883*4)+3] <= 1'b1;
                  spc883_inst_done         <= `ARIANE_CORE883.piton_pc_vld;
                  spc883_phy_pc_w          <= `ARIANE_CORE883.piton_pc;
                end
            end
    

            assign spc884_thread_id = 2'b00;
            assign spc884_rtl_pc = spc884_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(884*4)]   <= 1'b0;
                  active_thread[(884*4)+1] <= 1'b0;
                  active_thread[(884*4)+2] <= 1'b0;
                  active_thread[(884*4)+3] <= 1'b0;
                  spc884_inst_done         <= 0;
                  spc884_phy_pc_w          <= 0;
                end else begin
                  active_thread[(884*4)]   <= 1'b1;
                  active_thread[(884*4)+1] <= 1'b1;
                  active_thread[(884*4)+2] <= 1'b1;
                  active_thread[(884*4)+3] <= 1'b1;
                  spc884_inst_done         <= `ARIANE_CORE884.piton_pc_vld;
                  spc884_phy_pc_w          <= `ARIANE_CORE884.piton_pc;
                end
            end
    

            assign spc885_thread_id = 2'b00;
            assign spc885_rtl_pc = spc885_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(885*4)]   <= 1'b0;
                  active_thread[(885*4)+1] <= 1'b0;
                  active_thread[(885*4)+2] <= 1'b0;
                  active_thread[(885*4)+3] <= 1'b0;
                  spc885_inst_done         <= 0;
                  spc885_phy_pc_w          <= 0;
                end else begin
                  active_thread[(885*4)]   <= 1'b1;
                  active_thread[(885*4)+1] <= 1'b1;
                  active_thread[(885*4)+2] <= 1'b1;
                  active_thread[(885*4)+3] <= 1'b1;
                  spc885_inst_done         <= `ARIANE_CORE885.piton_pc_vld;
                  spc885_phy_pc_w          <= `ARIANE_CORE885.piton_pc;
                end
            end
    

            assign spc886_thread_id = 2'b00;
            assign spc886_rtl_pc = spc886_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(886*4)]   <= 1'b0;
                  active_thread[(886*4)+1] <= 1'b0;
                  active_thread[(886*4)+2] <= 1'b0;
                  active_thread[(886*4)+3] <= 1'b0;
                  spc886_inst_done         <= 0;
                  spc886_phy_pc_w          <= 0;
                end else begin
                  active_thread[(886*4)]   <= 1'b1;
                  active_thread[(886*4)+1] <= 1'b1;
                  active_thread[(886*4)+2] <= 1'b1;
                  active_thread[(886*4)+3] <= 1'b1;
                  spc886_inst_done         <= `ARIANE_CORE886.piton_pc_vld;
                  spc886_phy_pc_w          <= `ARIANE_CORE886.piton_pc;
                end
            end
    

            assign spc887_thread_id = 2'b00;
            assign spc887_rtl_pc = spc887_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(887*4)]   <= 1'b0;
                  active_thread[(887*4)+1] <= 1'b0;
                  active_thread[(887*4)+2] <= 1'b0;
                  active_thread[(887*4)+3] <= 1'b0;
                  spc887_inst_done         <= 0;
                  spc887_phy_pc_w          <= 0;
                end else begin
                  active_thread[(887*4)]   <= 1'b1;
                  active_thread[(887*4)+1] <= 1'b1;
                  active_thread[(887*4)+2] <= 1'b1;
                  active_thread[(887*4)+3] <= 1'b1;
                  spc887_inst_done         <= `ARIANE_CORE887.piton_pc_vld;
                  spc887_phy_pc_w          <= `ARIANE_CORE887.piton_pc;
                end
            end
    

            assign spc888_thread_id = 2'b00;
            assign spc888_rtl_pc = spc888_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(888*4)]   <= 1'b0;
                  active_thread[(888*4)+1] <= 1'b0;
                  active_thread[(888*4)+2] <= 1'b0;
                  active_thread[(888*4)+3] <= 1'b0;
                  spc888_inst_done         <= 0;
                  spc888_phy_pc_w          <= 0;
                end else begin
                  active_thread[(888*4)]   <= 1'b1;
                  active_thread[(888*4)+1] <= 1'b1;
                  active_thread[(888*4)+2] <= 1'b1;
                  active_thread[(888*4)+3] <= 1'b1;
                  spc888_inst_done         <= `ARIANE_CORE888.piton_pc_vld;
                  spc888_phy_pc_w          <= `ARIANE_CORE888.piton_pc;
                end
            end
    

            assign spc889_thread_id = 2'b00;
            assign spc889_rtl_pc = spc889_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(889*4)]   <= 1'b0;
                  active_thread[(889*4)+1] <= 1'b0;
                  active_thread[(889*4)+2] <= 1'b0;
                  active_thread[(889*4)+3] <= 1'b0;
                  spc889_inst_done         <= 0;
                  spc889_phy_pc_w          <= 0;
                end else begin
                  active_thread[(889*4)]   <= 1'b1;
                  active_thread[(889*4)+1] <= 1'b1;
                  active_thread[(889*4)+2] <= 1'b1;
                  active_thread[(889*4)+3] <= 1'b1;
                  spc889_inst_done         <= `ARIANE_CORE889.piton_pc_vld;
                  spc889_phy_pc_w          <= `ARIANE_CORE889.piton_pc;
                end
            end
    

            assign spc890_thread_id = 2'b00;
            assign spc890_rtl_pc = spc890_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(890*4)]   <= 1'b0;
                  active_thread[(890*4)+1] <= 1'b0;
                  active_thread[(890*4)+2] <= 1'b0;
                  active_thread[(890*4)+3] <= 1'b0;
                  spc890_inst_done         <= 0;
                  spc890_phy_pc_w          <= 0;
                end else begin
                  active_thread[(890*4)]   <= 1'b1;
                  active_thread[(890*4)+1] <= 1'b1;
                  active_thread[(890*4)+2] <= 1'b1;
                  active_thread[(890*4)+3] <= 1'b1;
                  spc890_inst_done         <= `ARIANE_CORE890.piton_pc_vld;
                  spc890_phy_pc_w          <= `ARIANE_CORE890.piton_pc;
                end
            end
    

            assign spc891_thread_id = 2'b00;
            assign spc891_rtl_pc = spc891_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(891*4)]   <= 1'b0;
                  active_thread[(891*4)+1] <= 1'b0;
                  active_thread[(891*4)+2] <= 1'b0;
                  active_thread[(891*4)+3] <= 1'b0;
                  spc891_inst_done         <= 0;
                  spc891_phy_pc_w          <= 0;
                end else begin
                  active_thread[(891*4)]   <= 1'b1;
                  active_thread[(891*4)+1] <= 1'b1;
                  active_thread[(891*4)+2] <= 1'b1;
                  active_thread[(891*4)+3] <= 1'b1;
                  spc891_inst_done         <= `ARIANE_CORE891.piton_pc_vld;
                  spc891_phy_pc_w          <= `ARIANE_CORE891.piton_pc;
                end
            end
    

            assign spc892_thread_id = 2'b00;
            assign spc892_rtl_pc = spc892_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(892*4)]   <= 1'b0;
                  active_thread[(892*4)+1] <= 1'b0;
                  active_thread[(892*4)+2] <= 1'b0;
                  active_thread[(892*4)+3] <= 1'b0;
                  spc892_inst_done         <= 0;
                  spc892_phy_pc_w          <= 0;
                end else begin
                  active_thread[(892*4)]   <= 1'b1;
                  active_thread[(892*4)+1] <= 1'b1;
                  active_thread[(892*4)+2] <= 1'b1;
                  active_thread[(892*4)+3] <= 1'b1;
                  spc892_inst_done         <= `ARIANE_CORE892.piton_pc_vld;
                  spc892_phy_pc_w          <= `ARIANE_CORE892.piton_pc;
                end
            end
    

            assign spc893_thread_id = 2'b00;
            assign spc893_rtl_pc = spc893_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(893*4)]   <= 1'b0;
                  active_thread[(893*4)+1] <= 1'b0;
                  active_thread[(893*4)+2] <= 1'b0;
                  active_thread[(893*4)+3] <= 1'b0;
                  spc893_inst_done         <= 0;
                  spc893_phy_pc_w          <= 0;
                end else begin
                  active_thread[(893*4)]   <= 1'b1;
                  active_thread[(893*4)+1] <= 1'b1;
                  active_thread[(893*4)+2] <= 1'b1;
                  active_thread[(893*4)+3] <= 1'b1;
                  spc893_inst_done         <= `ARIANE_CORE893.piton_pc_vld;
                  spc893_phy_pc_w          <= `ARIANE_CORE893.piton_pc;
                end
            end
    

            assign spc894_thread_id = 2'b00;
            assign spc894_rtl_pc = spc894_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(894*4)]   <= 1'b0;
                  active_thread[(894*4)+1] <= 1'b0;
                  active_thread[(894*4)+2] <= 1'b0;
                  active_thread[(894*4)+3] <= 1'b0;
                  spc894_inst_done         <= 0;
                  spc894_phy_pc_w          <= 0;
                end else begin
                  active_thread[(894*4)]   <= 1'b1;
                  active_thread[(894*4)+1] <= 1'b1;
                  active_thread[(894*4)+2] <= 1'b1;
                  active_thread[(894*4)+3] <= 1'b1;
                  spc894_inst_done         <= `ARIANE_CORE894.piton_pc_vld;
                  spc894_phy_pc_w          <= `ARIANE_CORE894.piton_pc;
                end
            end
    

            assign spc895_thread_id = 2'b00;
            assign spc895_rtl_pc = spc895_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(895*4)]   <= 1'b0;
                  active_thread[(895*4)+1] <= 1'b0;
                  active_thread[(895*4)+2] <= 1'b0;
                  active_thread[(895*4)+3] <= 1'b0;
                  spc895_inst_done         <= 0;
                  spc895_phy_pc_w          <= 0;
                end else begin
                  active_thread[(895*4)]   <= 1'b1;
                  active_thread[(895*4)+1] <= 1'b1;
                  active_thread[(895*4)+2] <= 1'b1;
                  active_thread[(895*4)+3] <= 1'b1;
                  spc895_inst_done         <= `ARIANE_CORE895.piton_pc_vld;
                  spc895_phy_pc_w          <= `ARIANE_CORE895.piton_pc;
                end
            end
    

            assign spc896_thread_id = 2'b00;
            assign spc896_rtl_pc = spc896_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(896*4)]   <= 1'b0;
                  active_thread[(896*4)+1] <= 1'b0;
                  active_thread[(896*4)+2] <= 1'b0;
                  active_thread[(896*4)+3] <= 1'b0;
                  spc896_inst_done         <= 0;
                  spc896_phy_pc_w          <= 0;
                end else begin
                  active_thread[(896*4)]   <= 1'b1;
                  active_thread[(896*4)+1] <= 1'b1;
                  active_thread[(896*4)+2] <= 1'b1;
                  active_thread[(896*4)+3] <= 1'b1;
                  spc896_inst_done         <= `ARIANE_CORE896.piton_pc_vld;
                  spc896_phy_pc_w          <= `ARIANE_CORE896.piton_pc;
                end
            end
    

            assign spc897_thread_id = 2'b00;
            assign spc897_rtl_pc = spc897_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(897*4)]   <= 1'b0;
                  active_thread[(897*4)+1] <= 1'b0;
                  active_thread[(897*4)+2] <= 1'b0;
                  active_thread[(897*4)+3] <= 1'b0;
                  spc897_inst_done         <= 0;
                  spc897_phy_pc_w          <= 0;
                end else begin
                  active_thread[(897*4)]   <= 1'b1;
                  active_thread[(897*4)+1] <= 1'b1;
                  active_thread[(897*4)+2] <= 1'b1;
                  active_thread[(897*4)+3] <= 1'b1;
                  spc897_inst_done         <= `ARIANE_CORE897.piton_pc_vld;
                  spc897_phy_pc_w          <= `ARIANE_CORE897.piton_pc;
                end
            end
    

            assign spc898_thread_id = 2'b00;
            assign spc898_rtl_pc = spc898_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(898*4)]   <= 1'b0;
                  active_thread[(898*4)+1] <= 1'b0;
                  active_thread[(898*4)+2] <= 1'b0;
                  active_thread[(898*4)+3] <= 1'b0;
                  spc898_inst_done         <= 0;
                  spc898_phy_pc_w          <= 0;
                end else begin
                  active_thread[(898*4)]   <= 1'b1;
                  active_thread[(898*4)+1] <= 1'b1;
                  active_thread[(898*4)+2] <= 1'b1;
                  active_thread[(898*4)+3] <= 1'b1;
                  spc898_inst_done         <= `ARIANE_CORE898.piton_pc_vld;
                  spc898_phy_pc_w          <= `ARIANE_CORE898.piton_pc;
                end
            end
    

            assign spc899_thread_id = 2'b00;
            assign spc899_rtl_pc = spc899_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(899*4)]   <= 1'b0;
                  active_thread[(899*4)+1] <= 1'b0;
                  active_thread[(899*4)+2] <= 1'b0;
                  active_thread[(899*4)+3] <= 1'b0;
                  spc899_inst_done         <= 0;
                  spc899_phy_pc_w          <= 0;
                end else begin
                  active_thread[(899*4)]   <= 1'b1;
                  active_thread[(899*4)+1] <= 1'b1;
                  active_thread[(899*4)+2] <= 1'b1;
                  active_thread[(899*4)+3] <= 1'b1;
                  spc899_inst_done         <= `ARIANE_CORE899.piton_pc_vld;
                  spc899_phy_pc_w          <= `ARIANE_CORE899.piton_pc;
                end
            end
    

            assign spc900_thread_id = 2'b00;
            assign spc900_rtl_pc = spc900_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(900*4)]   <= 1'b0;
                  active_thread[(900*4)+1] <= 1'b0;
                  active_thread[(900*4)+2] <= 1'b0;
                  active_thread[(900*4)+3] <= 1'b0;
                  spc900_inst_done         <= 0;
                  spc900_phy_pc_w          <= 0;
                end else begin
                  active_thread[(900*4)]   <= 1'b1;
                  active_thread[(900*4)+1] <= 1'b1;
                  active_thread[(900*4)+2] <= 1'b1;
                  active_thread[(900*4)+3] <= 1'b1;
                  spc900_inst_done         <= `ARIANE_CORE900.piton_pc_vld;
                  spc900_phy_pc_w          <= `ARIANE_CORE900.piton_pc;
                end
            end
    

            assign spc901_thread_id = 2'b00;
            assign spc901_rtl_pc = spc901_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(901*4)]   <= 1'b0;
                  active_thread[(901*4)+1] <= 1'b0;
                  active_thread[(901*4)+2] <= 1'b0;
                  active_thread[(901*4)+3] <= 1'b0;
                  spc901_inst_done         <= 0;
                  spc901_phy_pc_w          <= 0;
                end else begin
                  active_thread[(901*4)]   <= 1'b1;
                  active_thread[(901*4)+1] <= 1'b1;
                  active_thread[(901*4)+2] <= 1'b1;
                  active_thread[(901*4)+3] <= 1'b1;
                  spc901_inst_done         <= `ARIANE_CORE901.piton_pc_vld;
                  spc901_phy_pc_w          <= `ARIANE_CORE901.piton_pc;
                end
            end
    

            assign spc902_thread_id = 2'b00;
            assign spc902_rtl_pc = spc902_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(902*4)]   <= 1'b0;
                  active_thread[(902*4)+1] <= 1'b0;
                  active_thread[(902*4)+2] <= 1'b0;
                  active_thread[(902*4)+3] <= 1'b0;
                  spc902_inst_done         <= 0;
                  spc902_phy_pc_w          <= 0;
                end else begin
                  active_thread[(902*4)]   <= 1'b1;
                  active_thread[(902*4)+1] <= 1'b1;
                  active_thread[(902*4)+2] <= 1'b1;
                  active_thread[(902*4)+3] <= 1'b1;
                  spc902_inst_done         <= `ARIANE_CORE902.piton_pc_vld;
                  spc902_phy_pc_w          <= `ARIANE_CORE902.piton_pc;
                end
            end
    

            assign spc903_thread_id = 2'b00;
            assign spc903_rtl_pc = spc903_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(903*4)]   <= 1'b0;
                  active_thread[(903*4)+1] <= 1'b0;
                  active_thread[(903*4)+2] <= 1'b0;
                  active_thread[(903*4)+3] <= 1'b0;
                  spc903_inst_done         <= 0;
                  spc903_phy_pc_w          <= 0;
                end else begin
                  active_thread[(903*4)]   <= 1'b1;
                  active_thread[(903*4)+1] <= 1'b1;
                  active_thread[(903*4)+2] <= 1'b1;
                  active_thread[(903*4)+3] <= 1'b1;
                  spc903_inst_done         <= `ARIANE_CORE903.piton_pc_vld;
                  spc903_phy_pc_w          <= `ARIANE_CORE903.piton_pc;
                end
            end
    

            assign spc904_thread_id = 2'b00;
            assign spc904_rtl_pc = spc904_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(904*4)]   <= 1'b0;
                  active_thread[(904*4)+1] <= 1'b0;
                  active_thread[(904*4)+2] <= 1'b0;
                  active_thread[(904*4)+3] <= 1'b0;
                  spc904_inst_done         <= 0;
                  spc904_phy_pc_w          <= 0;
                end else begin
                  active_thread[(904*4)]   <= 1'b1;
                  active_thread[(904*4)+1] <= 1'b1;
                  active_thread[(904*4)+2] <= 1'b1;
                  active_thread[(904*4)+3] <= 1'b1;
                  spc904_inst_done         <= `ARIANE_CORE904.piton_pc_vld;
                  spc904_phy_pc_w          <= `ARIANE_CORE904.piton_pc;
                end
            end
    

            assign spc905_thread_id = 2'b00;
            assign spc905_rtl_pc = spc905_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(905*4)]   <= 1'b0;
                  active_thread[(905*4)+1] <= 1'b0;
                  active_thread[(905*4)+2] <= 1'b0;
                  active_thread[(905*4)+3] <= 1'b0;
                  spc905_inst_done         <= 0;
                  spc905_phy_pc_w          <= 0;
                end else begin
                  active_thread[(905*4)]   <= 1'b1;
                  active_thread[(905*4)+1] <= 1'b1;
                  active_thread[(905*4)+2] <= 1'b1;
                  active_thread[(905*4)+3] <= 1'b1;
                  spc905_inst_done         <= `ARIANE_CORE905.piton_pc_vld;
                  spc905_phy_pc_w          <= `ARIANE_CORE905.piton_pc;
                end
            end
    

            assign spc906_thread_id = 2'b00;
            assign spc906_rtl_pc = spc906_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(906*4)]   <= 1'b0;
                  active_thread[(906*4)+1] <= 1'b0;
                  active_thread[(906*4)+2] <= 1'b0;
                  active_thread[(906*4)+3] <= 1'b0;
                  spc906_inst_done         <= 0;
                  spc906_phy_pc_w          <= 0;
                end else begin
                  active_thread[(906*4)]   <= 1'b1;
                  active_thread[(906*4)+1] <= 1'b1;
                  active_thread[(906*4)+2] <= 1'b1;
                  active_thread[(906*4)+3] <= 1'b1;
                  spc906_inst_done         <= `ARIANE_CORE906.piton_pc_vld;
                  spc906_phy_pc_w          <= `ARIANE_CORE906.piton_pc;
                end
            end
    

            assign spc907_thread_id = 2'b00;
            assign spc907_rtl_pc = spc907_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(907*4)]   <= 1'b0;
                  active_thread[(907*4)+1] <= 1'b0;
                  active_thread[(907*4)+2] <= 1'b0;
                  active_thread[(907*4)+3] <= 1'b0;
                  spc907_inst_done         <= 0;
                  spc907_phy_pc_w          <= 0;
                end else begin
                  active_thread[(907*4)]   <= 1'b1;
                  active_thread[(907*4)+1] <= 1'b1;
                  active_thread[(907*4)+2] <= 1'b1;
                  active_thread[(907*4)+3] <= 1'b1;
                  spc907_inst_done         <= `ARIANE_CORE907.piton_pc_vld;
                  spc907_phy_pc_w          <= `ARIANE_CORE907.piton_pc;
                end
            end
    

            assign spc908_thread_id = 2'b00;
            assign spc908_rtl_pc = spc908_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(908*4)]   <= 1'b0;
                  active_thread[(908*4)+1] <= 1'b0;
                  active_thread[(908*4)+2] <= 1'b0;
                  active_thread[(908*4)+3] <= 1'b0;
                  spc908_inst_done         <= 0;
                  spc908_phy_pc_w          <= 0;
                end else begin
                  active_thread[(908*4)]   <= 1'b1;
                  active_thread[(908*4)+1] <= 1'b1;
                  active_thread[(908*4)+2] <= 1'b1;
                  active_thread[(908*4)+3] <= 1'b1;
                  spc908_inst_done         <= `ARIANE_CORE908.piton_pc_vld;
                  spc908_phy_pc_w          <= `ARIANE_CORE908.piton_pc;
                end
            end
    

            assign spc909_thread_id = 2'b00;
            assign spc909_rtl_pc = spc909_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(909*4)]   <= 1'b0;
                  active_thread[(909*4)+1] <= 1'b0;
                  active_thread[(909*4)+2] <= 1'b0;
                  active_thread[(909*4)+3] <= 1'b0;
                  spc909_inst_done         <= 0;
                  spc909_phy_pc_w          <= 0;
                end else begin
                  active_thread[(909*4)]   <= 1'b1;
                  active_thread[(909*4)+1] <= 1'b1;
                  active_thread[(909*4)+2] <= 1'b1;
                  active_thread[(909*4)+3] <= 1'b1;
                  spc909_inst_done         <= `ARIANE_CORE909.piton_pc_vld;
                  spc909_phy_pc_w          <= `ARIANE_CORE909.piton_pc;
                end
            end
    

            assign spc910_thread_id = 2'b00;
            assign spc910_rtl_pc = spc910_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(910*4)]   <= 1'b0;
                  active_thread[(910*4)+1] <= 1'b0;
                  active_thread[(910*4)+2] <= 1'b0;
                  active_thread[(910*4)+3] <= 1'b0;
                  spc910_inst_done         <= 0;
                  spc910_phy_pc_w          <= 0;
                end else begin
                  active_thread[(910*4)]   <= 1'b1;
                  active_thread[(910*4)+1] <= 1'b1;
                  active_thread[(910*4)+2] <= 1'b1;
                  active_thread[(910*4)+3] <= 1'b1;
                  spc910_inst_done         <= `ARIANE_CORE910.piton_pc_vld;
                  spc910_phy_pc_w          <= `ARIANE_CORE910.piton_pc;
                end
            end
    

            assign spc911_thread_id = 2'b00;
            assign spc911_rtl_pc = spc911_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(911*4)]   <= 1'b0;
                  active_thread[(911*4)+1] <= 1'b0;
                  active_thread[(911*4)+2] <= 1'b0;
                  active_thread[(911*4)+3] <= 1'b0;
                  spc911_inst_done         <= 0;
                  spc911_phy_pc_w          <= 0;
                end else begin
                  active_thread[(911*4)]   <= 1'b1;
                  active_thread[(911*4)+1] <= 1'b1;
                  active_thread[(911*4)+2] <= 1'b1;
                  active_thread[(911*4)+3] <= 1'b1;
                  spc911_inst_done         <= `ARIANE_CORE911.piton_pc_vld;
                  spc911_phy_pc_w          <= `ARIANE_CORE911.piton_pc;
                end
            end
    

            assign spc912_thread_id = 2'b00;
            assign spc912_rtl_pc = spc912_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(912*4)]   <= 1'b0;
                  active_thread[(912*4)+1] <= 1'b0;
                  active_thread[(912*4)+2] <= 1'b0;
                  active_thread[(912*4)+3] <= 1'b0;
                  spc912_inst_done         <= 0;
                  spc912_phy_pc_w          <= 0;
                end else begin
                  active_thread[(912*4)]   <= 1'b1;
                  active_thread[(912*4)+1] <= 1'b1;
                  active_thread[(912*4)+2] <= 1'b1;
                  active_thread[(912*4)+3] <= 1'b1;
                  spc912_inst_done         <= `ARIANE_CORE912.piton_pc_vld;
                  spc912_phy_pc_w          <= `ARIANE_CORE912.piton_pc;
                end
            end
    

            assign spc913_thread_id = 2'b00;
            assign spc913_rtl_pc = spc913_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(913*4)]   <= 1'b0;
                  active_thread[(913*4)+1] <= 1'b0;
                  active_thread[(913*4)+2] <= 1'b0;
                  active_thread[(913*4)+3] <= 1'b0;
                  spc913_inst_done         <= 0;
                  spc913_phy_pc_w          <= 0;
                end else begin
                  active_thread[(913*4)]   <= 1'b1;
                  active_thread[(913*4)+1] <= 1'b1;
                  active_thread[(913*4)+2] <= 1'b1;
                  active_thread[(913*4)+3] <= 1'b1;
                  spc913_inst_done         <= `ARIANE_CORE913.piton_pc_vld;
                  spc913_phy_pc_w          <= `ARIANE_CORE913.piton_pc;
                end
            end
    

            assign spc914_thread_id = 2'b00;
            assign spc914_rtl_pc = spc914_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(914*4)]   <= 1'b0;
                  active_thread[(914*4)+1] <= 1'b0;
                  active_thread[(914*4)+2] <= 1'b0;
                  active_thread[(914*4)+3] <= 1'b0;
                  spc914_inst_done         <= 0;
                  spc914_phy_pc_w          <= 0;
                end else begin
                  active_thread[(914*4)]   <= 1'b1;
                  active_thread[(914*4)+1] <= 1'b1;
                  active_thread[(914*4)+2] <= 1'b1;
                  active_thread[(914*4)+3] <= 1'b1;
                  spc914_inst_done         <= `ARIANE_CORE914.piton_pc_vld;
                  spc914_phy_pc_w          <= `ARIANE_CORE914.piton_pc;
                end
            end
    

            assign spc915_thread_id = 2'b00;
            assign spc915_rtl_pc = spc915_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(915*4)]   <= 1'b0;
                  active_thread[(915*4)+1] <= 1'b0;
                  active_thread[(915*4)+2] <= 1'b0;
                  active_thread[(915*4)+3] <= 1'b0;
                  spc915_inst_done         <= 0;
                  spc915_phy_pc_w          <= 0;
                end else begin
                  active_thread[(915*4)]   <= 1'b1;
                  active_thread[(915*4)+1] <= 1'b1;
                  active_thread[(915*4)+2] <= 1'b1;
                  active_thread[(915*4)+3] <= 1'b1;
                  spc915_inst_done         <= `ARIANE_CORE915.piton_pc_vld;
                  spc915_phy_pc_w          <= `ARIANE_CORE915.piton_pc;
                end
            end
    

            assign spc916_thread_id = 2'b00;
            assign spc916_rtl_pc = spc916_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(916*4)]   <= 1'b0;
                  active_thread[(916*4)+1] <= 1'b0;
                  active_thread[(916*4)+2] <= 1'b0;
                  active_thread[(916*4)+3] <= 1'b0;
                  spc916_inst_done         <= 0;
                  spc916_phy_pc_w          <= 0;
                end else begin
                  active_thread[(916*4)]   <= 1'b1;
                  active_thread[(916*4)+1] <= 1'b1;
                  active_thread[(916*4)+2] <= 1'b1;
                  active_thread[(916*4)+3] <= 1'b1;
                  spc916_inst_done         <= `ARIANE_CORE916.piton_pc_vld;
                  spc916_phy_pc_w          <= `ARIANE_CORE916.piton_pc;
                end
            end
    

            assign spc917_thread_id = 2'b00;
            assign spc917_rtl_pc = spc917_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(917*4)]   <= 1'b0;
                  active_thread[(917*4)+1] <= 1'b0;
                  active_thread[(917*4)+2] <= 1'b0;
                  active_thread[(917*4)+3] <= 1'b0;
                  spc917_inst_done         <= 0;
                  spc917_phy_pc_w          <= 0;
                end else begin
                  active_thread[(917*4)]   <= 1'b1;
                  active_thread[(917*4)+1] <= 1'b1;
                  active_thread[(917*4)+2] <= 1'b1;
                  active_thread[(917*4)+3] <= 1'b1;
                  spc917_inst_done         <= `ARIANE_CORE917.piton_pc_vld;
                  spc917_phy_pc_w          <= `ARIANE_CORE917.piton_pc;
                end
            end
    

            assign spc918_thread_id = 2'b00;
            assign spc918_rtl_pc = spc918_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(918*4)]   <= 1'b0;
                  active_thread[(918*4)+1] <= 1'b0;
                  active_thread[(918*4)+2] <= 1'b0;
                  active_thread[(918*4)+3] <= 1'b0;
                  spc918_inst_done         <= 0;
                  spc918_phy_pc_w          <= 0;
                end else begin
                  active_thread[(918*4)]   <= 1'b1;
                  active_thread[(918*4)+1] <= 1'b1;
                  active_thread[(918*4)+2] <= 1'b1;
                  active_thread[(918*4)+3] <= 1'b1;
                  spc918_inst_done         <= `ARIANE_CORE918.piton_pc_vld;
                  spc918_phy_pc_w          <= `ARIANE_CORE918.piton_pc;
                end
            end
    

            assign spc919_thread_id = 2'b00;
            assign spc919_rtl_pc = spc919_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(919*4)]   <= 1'b0;
                  active_thread[(919*4)+1] <= 1'b0;
                  active_thread[(919*4)+2] <= 1'b0;
                  active_thread[(919*4)+3] <= 1'b0;
                  spc919_inst_done         <= 0;
                  spc919_phy_pc_w          <= 0;
                end else begin
                  active_thread[(919*4)]   <= 1'b1;
                  active_thread[(919*4)+1] <= 1'b1;
                  active_thread[(919*4)+2] <= 1'b1;
                  active_thread[(919*4)+3] <= 1'b1;
                  spc919_inst_done         <= `ARIANE_CORE919.piton_pc_vld;
                  spc919_phy_pc_w          <= `ARIANE_CORE919.piton_pc;
                end
            end
    

            assign spc920_thread_id = 2'b00;
            assign spc920_rtl_pc = spc920_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(920*4)]   <= 1'b0;
                  active_thread[(920*4)+1] <= 1'b0;
                  active_thread[(920*4)+2] <= 1'b0;
                  active_thread[(920*4)+3] <= 1'b0;
                  spc920_inst_done         <= 0;
                  spc920_phy_pc_w          <= 0;
                end else begin
                  active_thread[(920*4)]   <= 1'b1;
                  active_thread[(920*4)+1] <= 1'b1;
                  active_thread[(920*4)+2] <= 1'b1;
                  active_thread[(920*4)+3] <= 1'b1;
                  spc920_inst_done         <= `ARIANE_CORE920.piton_pc_vld;
                  spc920_phy_pc_w          <= `ARIANE_CORE920.piton_pc;
                end
            end
    

            assign spc921_thread_id = 2'b00;
            assign spc921_rtl_pc = spc921_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(921*4)]   <= 1'b0;
                  active_thread[(921*4)+1] <= 1'b0;
                  active_thread[(921*4)+2] <= 1'b0;
                  active_thread[(921*4)+3] <= 1'b0;
                  spc921_inst_done         <= 0;
                  spc921_phy_pc_w          <= 0;
                end else begin
                  active_thread[(921*4)]   <= 1'b1;
                  active_thread[(921*4)+1] <= 1'b1;
                  active_thread[(921*4)+2] <= 1'b1;
                  active_thread[(921*4)+3] <= 1'b1;
                  spc921_inst_done         <= `ARIANE_CORE921.piton_pc_vld;
                  spc921_phy_pc_w          <= `ARIANE_CORE921.piton_pc;
                end
            end
    

            assign spc922_thread_id = 2'b00;
            assign spc922_rtl_pc = spc922_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(922*4)]   <= 1'b0;
                  active_thread[(922*4)+1] <= 1'b0;
                  active_thread[(922*4)+2] <= 1'b0;
                  active_thread[(922*4)+3] <= 1'b0;
                  spc922_inst_done         <= 0;
                  spc922_phy_pc_w          <= 0;
                end else begin
                  active_thread[(922*4)]   <= 1'b1;
                  active_thread[(922*4)+1] <= 1'b1;
                  active_thread[(922*4)+2] <= 1'b1;
                  active_thread[(922*4)+3] <= 1'b1;
                  spc922_inst_done         <= `ARIANE_CORE922.piton_pc_vld;
                  spc922_phy_pc_w          <= `ARIANE_CORE922.piton_pc;
                end
            end
    

            assign spc923_thread_id = 2'b00;
            assign spc923_rtl_pc = spc923_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(923*4)]   <= 1'b0;
                  active_thread[(923*4)+1] <= 1'b0;
                  active_thread[(923*4)+2] <= 1'b0;
                  active_thread[(923*4)+3] <= 1'b0;
                  spc923_inst_done         <= 0;
                  spc923_phy_pc_w          <= 0;
                end else begin
                  active_thread[(923*4)]   <= 1'b1;
                  active_thread[(923*4)+1] <= 1'b1;
                  active_thread[(923*4)+2] <= 1'b1;
                  active_thread[(923*4)+3] <= 1'b1;
                  spc923_inst_done         <= `ARIANE_CORE923.piton_pc_vld;
                  spc923_phy_pc_w          <= `ARIANE_CORE923.piton_pc;
                end
            end
    

            assign spc924_thread_id = 2'b00;
            assign spc924_rtl_pc = spc924_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(924*4)]   <= 1'b0;
                  active_thread[(924*4)+1] <= 1'b0;
                  active_thread[(924*4)+2] <= 1'b0;
                  active_thread[(924*4)+3] <= 1'b0;
                  spc924_inst_done         <= 0;
                  spc924_phy_pc_w          <= 0;
                end else begin
                  active_thread[(924*4)]   <= 1'b1;
                  active_thread[(924*4)+1] <= 1'b1;
                  active_thread[(924*4)+2] <= 1'b1;
                  active_thread[(924*4)+3] <= 1'b1;
                  spc924_inst_done         <= `ARIANE_CORE924.piton_pc_vld;
                  spc924_phy_pc_w          <= `ARIANE_CORE924.piton_pc;
                end
            end
    

            assign spc925_thread_id = 2'b00;
            assign spc925_rtl_pc = spc925_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(925*4)]   <= 1'b0;
                  active_thread[(925*4)+1] <= 1'b0;
                  active_thread[(925*4)+2] <= 1'b0;
                  active_thread[(925*4)+3] <= 1'b0;
                  spc925_inst_done         <= 0;
                  spc925_phy_pc_w          <= 0;
                end else begin
                  active_thread[(925*4)]   <= 1'b1;
                  active_thread[(925*4)+1] <= 1'b1;
                  active_thread[(925*4)+2] <= 1'b1;
                  active_thread[(925*4)+3] <= 1'b1;
                  spc925_inst_done         <= `ARIANE_CORE925.piton_pc_vld;
                  spc925_phy_pc_w          <= `ARIANE_CORE925.piton_pc;
                end
            end
    

            assign spc926_thread_id = 2'b00;
            assign spc926_rtl_pc = spc926_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(926*4)]   <= 1'b0;
                  active_thread[(926*4)+1] <= 1'b0;
                  active_thread[(926*4)+2] <= 1'b0;
                  active_thread[(926*4)+3] <= 1'b0;
                  spc926_inst_done         <= 0;
                  spc926_phy_pc_w          <= 0;
                end else begin
                  active_thread[(926*4)]   <= 1'b1;
                  active_thread[(926*4)+1] <= 1'b1;
                  active_thread[(926*4)+2] <= 1'b1;
                  active_thread[(926*4)+3] <= 1'b1;
                  spc926_inst_done         <= `ARIANE_CORE926.piton_pc_vld;
                  spc926_phy_pc_w          <= `ARIANE_CORE926.piton_pc;
                end
            end
    

            assign spc927_thread_id = 2'b00;
            assign spc927_rtl_pc = spc927_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(927*4)]   <= 1'b0;
                  active_thread[(927*4)+1] <= 1'b0;
                  active_thread[(927*4)+2] <= 1'b0;
                  active_thread[(927*4)+3] <= 1'b0;
                  spc927_inst_done         <= 0;
                  spc927_phy_pc_w          <= 0;
                end else begin
                  active_thread[(927*4)]   <= 1'b1;
                  active_thread[(927*4)+1] <= 1'b1;
                  active_thread[(927*4)+2] <= 1'b1;
                  active_thread[(927*4)+3] <= 1'b1;
                  spc927_inst_done         <= `ARIANE_CORE927.piton_pc_vld;
                  spc927_phy_pc_w          <= `ARIANE_CORE927.piton_pc;
                end
            end
    

            assign spc928_thread_id = 2'b00;
            assign spc928_rtl_pc = spc928_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(928*4)]   <= 1'b0;
                  active_thread[(928*4)+1] <= 1'b0;
                  active_thread[(928*4)+2] <= 1'b0;
                  active_thread[(928*4)+3] <= 1'b0;
                  spc928_inst_done         <= 0;
                  spc928_phy_pc_w          <= 0;
                end else begin
                  active_thread[(928*4)]   <= 1'b1;
                  active_thread[(928*4)+1] <= 1'b1;
                  active_thread[(928*4)+2] <= 1'b1;
                  active_thread[(928*4)+3] <= 1'b1;
                  spc928_inst_done         <= `ARIANE_CORE928.piton_pc_vld;
                  spc928_phy_pc_w          <= `ARIANE_CORE928.piton_pc;
                end
            end
    

            assign spc929_thread_id = 2'b00;
            assign spc929_rtl_pc = spc929_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(929*4)]   <= 1'b0;
                  active_thread[(929*4)+1] <= 1'b0;
                  active_thread[(929*4)+2] <= 1'b0;
                  active_thread[(929*4)+3] <= 1'b0;
                  spc929_inst_done         <= 0;
                  spc929_phy_pc_w          <= 0;
                end else begin
                  active_thread[(929*4)]   <= 1'b1;
                  active_thread[(929*4)+1] <= 1'b1;
                  active_thread[(929*4)+2] <= 1'b1;
                  active_thread[(929*4)+3] <= 1'b1;
                  spc929_inst_done         <= `ARIANE_CORE929.piton_pc_vld;
                  spc929_phy_pc_w          <= `ARIANE_CORE929.piton_pc;
                end
            end
    

            assign spc930_thread_id = 2'b00;
            assign spc930_rtl_pc = spc930_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(930*4)]   <= 1'b0;
                  active_thread[(930*4)+1] <= 1'b0;
                  active_thread[(930*4)+2] <= 1'b0;
                  active_thread[(930*4)+3] <= 1'b0;
                  spc930_inst_done         <= 0;
                  spc930_phy_pc_w          <= 0;
                end else begin
                  active_thread[(930*4)]   <= 1'b1;
                  active_thread[(930*4)+1] <= 1'b1;
                  active_thread[(930*4)+2] <= 1'b1;
                  active_thread[(930*4)+3] <= 1'b1;
                  spc930_inst_done         <= `ARIANE_CORE930.piton_pc_vld;
                  spc930_phy_pc_w          <= `ARIANE_CORE930.piton_pc;
                end
            end
    

            assign spc931_thread_id = 2'b00;
            assign spc931_rtl_pc = spc931_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(931*4)]   <= 1'b0;
                  active_thread[(931*4)+1] <= 1'b0;
                  active_thread[(931*4)+2] <= 1'b0;
                  active_thread[(931*4)+3] <= 1'b0;
                  spc931_inst_done         <= 0;
                  spc931_phy_pc_w          <= 0;
                end else begin
                  active_thread[(931*4)]   <= 1'b1;
                  active_thread[(931*4)+1] <= 1'b1;
                  active_thread[(931*4)+2] <= 1'b1;
                  active_thread[(931*4)+3] <= 1'b1;
                  spc931_inst_done         <= `ARIANE_CORE931.piton_pc_vld;
                  spc931_phy_pc_w          <= `ARIANE_CORE931.piton_pc;
                end
            end
    

            assign spc932_thread_id = 2'b00;
            assign spc932_rtl_pc = spc932_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(932*4)]   <= 1'b0;
                  active_thread[(932*4)+1] <= 1'b0;
                  active_thread[(932*4)+2] <= 1'b0;
                  active_thread[(932*4)+3] <= 1'b0;
                  spc932_inst_done         <= 0;
                  spc932_phy_pc_w          <= 0;
                end else begin
                  active_thread[(932*4)]   <= 1'b1;
                  active_thread[(932*4)+1] <= 1'b1;
                  active_thread[(932*4)+2] <= 1'b1;
                  active_thread[(932*4)+3] <= 1'b1;
                  spc932_inst_done         <= `ARIANE_CORE932.piton_pc_vld;
                  spc932_phy_pc_w          <= `ARIANE_CORE932.piton_pc;
                end
            end
    

            assign spc933_thread_id = 2'b00;
            assign spc933_rtl_pc = spc933_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(933*4)]   <= 1'b0;
                  active_thread[(933*4)+1] <= 1'b0;
                  active_thread[(933*4)+2] <= 1'b0;
                  active_thread[(933*4)+3] <= 1'b0;
                  spc933_inst_done         <= 0;
                  spc933_phy_pc_w          <= 0;
                end else begin
                  active_thread[(933*4)]   <= 1'b1;
                  active_thread[(933*4)+1] <= 1'b1;
                  active_thread[(933*4)+2] <= 1'b1;
                  active_thread[(933*4)+3] <= 1'b1;
                  spc933_inst_done         <= `ARIANE_CORE933.piton_pc_vld;
                  spc933_phy_pc_w          <= `ARIANE_CORE933.piton_pc;
                end
            end
    

            assign spc934_thread_id = 2'b00;
            assign spc934_rtl_pc = spc934_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(934*4)]   <= 1'b0;
                  active_thread[(934*4)+1] <= 1'b0;
                  active_thread[(934*4)+2] <= 1'b0;
                  active_thread[(934*4)+3] <= 1'b0;
                  spc934_inst_done         <= 0;
                  spc934_phy_pc_w          <= 0;
                end else begin
                  active_thread[(934*4)]   <= 1'b1;
                  active_thread[(934*4)+1] <= 1'b1;
                  active_thread[(934*4)+2] <= 1'b1;
                  active_thread[(934*4)+3] <= 1'b1;
                  spc934_inst_done         <= `ARIANE_CORE934.piton_pc_vld;
                  spc934_phy_pc_w          <= `ARIANE_CORE934.piton_pc;
                end
            end
    

            assign spc935_thread_id = 2'b00;
            assign spc935_rtl_pc = spc935_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(935*4)]   <= 1'b0;
                  active_thread[(935*4)+1] <= 1'b0;
                  active_thread[(935*4)+2] <= 1'b0;
                  active_thread[(935*4)+3] <= 1'b0;
                  spc935_inst_done         <= 0;
                  spc935_phy_pc_w          <= 0;
                end else begin
                  active_thread[(935*4)]   <= 1'b1;
                  active_thread[(935*4)+1] <= 1'b1;
                  active_thread[(935*4)+2] <= 1'b1;
                  active_thread[(935*4)+3] <= 1'b1;
                  spc935_inst_done         <= `ARIANE_CORE935.piton_pc_vld;
                  spc935_phy_pc_w          <= `ARIANE_CORE935.piton_pc;
                end
            end
    

            assign spc936_thread_id = 2'b00;
            assign spc936_rtl_pc = spc936_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(936*4)]   <= 1'b0;
                  active_thread[(936*4)+1] <= 1'b0;
                  active_thread[(936*4)+2] <= 1'b0;
                  active_thread[(936*4)+3] <= 1'b0;
                  spc936_inst_done         <= 0;
                  spc936_phy_pc_w          <= 0;
                end else begin
                  active_thread[(936*4)]   <= 1'b1;
                  active_thread[(936*4)+1] <= 1'b1;
                  active_thread[(936*4)+2] <= 1'b1;
                  active_thread[(936*4)+3] <= 1'b1;
                  spc936_inst_done         <= `ARIANE_CORE936.piton_pc_vld;
                  spc936_phy_pc_w          <= `ARIANE_CORE936.piton_pc;
                end
            end
    

            assign spc937_thread_id = 2'b00;
            assign spc937_rtl_pc = spc937_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(937*4)]   <= 1'b0;
                  active_thread[(937*4)+1] <= 1'b0;
                  active_thread[(937*4)+2] <= 1'b0;
                  active_thread[(937*4)+3] <= 1'b0;
                  spc937_inst_done         <= 0;
                  spc937_phy_pc_w          <= 0;
                end else begin
                  active_thread[(937*4)]   <= 1'b1;
                  active_thread[(937*4)+1] <= 1'b1;
                  active_thread[(937*4)+2] <= 1'b1;
                  active_thread[(937*4)+3] <= 1'b1;
                  spc937_inst_done         <= `ARIANE_CORE937.piton_pc_vld;
                  spc937_phy_pc_w          <= `ARIANE_CORE937.piton_pc;
                end
            end
    

            assign spc938_thread_id = 2'b00;
            assign spc938_rtl_pc = spc938_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(938*4)]   <= 1'b0;
                  active_thread[(938*4)+1] <= 1'b0;
                  active_thread[(938*4)+2] <= 1'b0;
                  active_thread[(938*4)+3] <= 1'b0;
                  spc938_inst_done         <= 0;
                  spc938_phy_pc_w          <= 0;
                end else begin
                  active_thread[(938*4)]   <= 1'b1;
                  active_thread[(938*4)+1] <= 1'b1;
                  active_thread[(938*4)+2] <= 1'b1;
                  active_thread[(938*4)+3] <= 1'b1;
                  spc938_inst_done         <= `ARIANE_CORE938.piton_pc_vld;
                  spc938_phy_pc_w          <= `ARIANE_CORE938.piton_pc;
                end
            end
    

            assign spc939_thread_id = 2'b00;
            assign spc939_rtl_pc = spc939_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(939*4)]   <= 1'b0;
                  active_thread[(939*4)+1] <= 1'b0;
                  active_thread[(939*4)+2] <= 1'b0;
                  active_thread[(939*4)+3] <= 1'b0;
                  spc939_inst_done         <= 0;
                  spc939_phy_pc_w          <= 0;
                end else begin
                  active_thread[(939*4)]   <= 1'b1;
                  active_thread[(939*4)+1] <= 1'b1;
                  active_thread[(939*4)+2] <= 1'b1;
                  active_thread[(939*4)+3] <= 1'b1;
                  spc939_inst_done         <= `ARIANE_CORE939.piton_pc_vld;
                  spc939_phy_pc_w          <= `ARIANE_CORE939.piton_pc;
                end
            end
    

            assign spc940_thread_id = 2'b00;
            assign spc940_rtl_pc = spc940_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(940*4)]   <= 1'b0;
                  active_thread[(940*4)+1] <= 1'b0;
                  active_thread[(940*4)+2] <= 1'b0;
                  active_thread[(940*4)+3] <= 1'b0;
                  spc940_inst_done         <= 0;
                  spc940_phy_pc_w          <= 0;
                end else begin
                  active_thread[(940*4)]   <= 1'b1;
                  active_thread[(940*4)+1] <= 1'b1;
                  active_thread[(940*4)+2] <= 1'b1;
                  active_thread[(940*4)+3] <= 1'b1;
                  spc940_inst_done         <= `ARIANE_CORE940.piton_pc_vld;
                  spc940_phy_pc_w          <= `ARIANE_CORE940.piton_pc;
                end
            end
    

            assign spc941_thread_id = 2'b00;
            assign spc941_rtl_pc = spc941_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(941*4)]   <= 1'b0;
                  active_thread[(941*4)+1] <= 1'b0;
                  active_thread[(941*4)+2] <= 1'b0;
                  active_thread[(941*4)+3] <= 1'b0;
                  spc941_inst_done         <= 0;
                  spc941_phy_pc_w          <= 0;
                end else begin
                  active_thread[(941*4)]   <= 1'b1;
                  active_thread[(941*4)+1] <= 1'b1;
                  active_thread[(941*4)+2] <= 1'b1;
                  active_thread[(941*4)+3] <= 1'b1;
                  spc941_inst_done         <= `ARIANE_CORE941.piton_pc_vld;
                  spc941_phy_pc_w          <= `ARIANE_CORE941.piton_pc;
                end
            end
    

            assign spc942_thread_id = 2'b00;
            assign spc942_rtl_pc = spc942_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(942*4)]   <= 1'b0;
                  active_thread[(942*4)+1] <= 1'b0;
                  active_thread[(942*4)+2] <= 1'b0;
                  active_thread[(942*4)+3] <= 1'b0;
                  spc942_inst_done         <= 0;
                  spc942_phy_pc_w          <= 0;
                end else begin
                  active_thread[(942*4)]   <= 1'b1;
                  active_thread[(942*4)+1] <= 1'b1;
                  active_thread[(942*4)+2] <= 1'b1;
                  active_thread[(942*4)+3] <= 1'b1;
                  spc942_inst_done         <= `ARIANE_CORE942.piton_pc_vld;
                  spc942_phy_pc_w          <= `ARIANE_CORE942.piton_pc;
                end
            end
    

            assign spc943_thread_id = 2'b00;
            assign spc943_rtl_pc = spc943_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(943*4)]   <= 1'b0;
                  active_thread[(943*4)+1] <= 1'b0;
                  active_thread[(943*4)+2] <= 1'b0;
                  active_thread[(943*4)+3] <= 1'b0;
                  spc943_inst_done         <= 0;
                  spc943_phy_pc_w          <= 0;
                end else begin
                  active_thread[(943*4)]   <= 1'b1;
                  active_thread[(943*4)+1] <= 1'b1;
                  active_thread[(943*4)+2] <= 1'b1;
                  active_thread[(943*4)+3] <= 1'b1;
                  spc943_inst_done         <= `ARIANE_CORE943.piton_pc_vld;
                  spc943_phy_pc_w          <= `ARIANE_CORE943.piton_pc;
                end
            end
    

            assign spc944_thread_id = 2'b00;
            assign spc944_rtl_pc = spc944_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(944*4)]   <= 1'b0;
                  active_thread[(944*4)+1] <= 1'b0;
                  active_thread[(944*4)+2] <= 1'b0;
                  active_thread[(944*4)+3] <= 1'b0;
                  spc944_inst_done         <= 0;
                  spc944_phy_pc_w          <= 0;
                end else begin
                  active_thread[(944*4)]   <= 1'b1;
                  active_thread[(944*4)+1] <= 1'b1;
                  active_thread[(944*4)+2] <= 1'b1;
                  active_thread[(944*4)+3] <= 1'b1;
                  spc944_inst_done         <= `ARIANE_CORE944.piton_pc_vld;
                  spc944_phy_pc_w          <= `ARIANE_CORE944.piton_pc;
                end
            end
    

            assign spc945_thread_id = 2'b00;
            assign spc945_rtl_pc = spc945_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(945*4)]   <= 1'b0;
                  active_thread[(945*4)+1] <= 1'b0;
                  active_thread[(945*4)+2] <= 1'b0;
                  active_thread[(945*4)+3] <= 1'b0;
                  spc945_inst_done         <= 0;
                  spc945_phy_pc_w          <= 0;
                end else begin
                  active_thread[(945*4)]   <= 1'b1;
                  active_thread[(945*4)+1] <= 1'b1;
                  active_thread[(945*4)+2] <= 1'b1;
                  active_thread[(945*4)+3] <= 1'b1;
                  spc945_inst_done         <= `ARIANE_CORE945.piton_pc_vld;
                  spc945_phy_pc_w          <= `ARIANE_CORE945.piton_pc;
                end
            end
    

            assign spc946_thread_id = 2'b00;
            assign spc946_rtl_pc = spc946_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(946*4)]   <= 1'b0;
                  active_thread[(946*4)+1] <= 1'b0;
                  active_thread[(946*4)+2] <= 1'b0;
                  active_thread[(946*4)+3] <= 1'b0;
                  spc946_inst_done         <= 0;
                  spc946_phy_pc_w          <= 0;
                end else begin
                  active_thread[(946*4)]   <= 1'b1;
                  active_thread[(946*4)+1] <= 1'b1;
                  active_thread[(946*4)+2] <= 1'b1;
                  active_thread[(946*4)+3] <= 1'b1;
                  spc946_inst_done         <= `ARIANE_CORE946.piton_pc_vld;
                  spc946_phy_pc_w          <= `ARIANE_CORE946.piton_pc;
                end
            end
    

            assign spc947_thread_id = 2'b00;
            assign spc947_rtl_pc = spc947_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(947*4)]   <= 1'b0;
                  active_thread[(947*4)+1] <= 1'b0;
                  active_thread[(947*4)+2] <= 1'b0;
                  active_thread[(947*4)+3] <= 1'b0;
                  spc947_inst_done         <= 0;
                  spc947_phy_pc_w          <= 0;
                end else begin
                  active_thread[(947*4)]   <= 1'b1;
                  active_thread[(947*4)+1] <= 1'b1;
                  active_thread[(947*4)+2] <= 1'b1;
                  active_thread[(947*4)+3] <= 1'b1;
                  spc947_inst_done         <= `ARIANE_CORE947.piton_pc_vld;
                  spc947_phy_pc_w          <= `ARIANE_CORE947.piton_pc;
                end
            end
    

            assign spc948_thread_id = 2'b00;
            assign spc948_rtl_pc = spc948_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(948*4)]   <= 1'b0;
                  active_thread[(948*4)+1] <= 1'b0;
                  active_thread[(948*4)+2] <= 1'b0;
                  active_thread[(948*4)+3] <= 1'b0;
                  spc948_inst_done         <= 0;
                  spc948_phy_pc_w          <= 0;
                end else begin
                  active_thread[(948*4)]   <= 1'b1;
                  active_thread[(948*4)+1] <= 1'b1;
                  active_thread[(948*4)+2] <= 1'b1;
                  active_thread[(948*4)+3] <= 1'b1;
                  spc948_inst_done         <= `ARIANE_CORE948.piton_pc_vld;
                  spc948_phy_pc_w          <= `ARIANE_CORE948.piton_pc;
                end
            end
    

            assign spc949_thread_id = 2'b00;
            assign spc949_rtl_pc = spc949_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(949*4)]   <= 1'b0;
                  active_thread[(949*4)+1] <= 1'b0;
                  active_thread[(949*4)+2] <= 1'b0;
                  active_thread[(949*4)+3] <= 1'b0;
                  spc949_inst_done         <= 0;
                  spc949_phy_pc_w          <= 0;
                end else begin
                  active_thread[(949*4)]   <= 1'b1;
                  active_thread[(949*4)+1] <= 1'b1;
                  active_thread[(949*4)+2] <= 1'b1;
                  active_thread[(949*4)+3] <= 1'b1;
                  spc949_inst_done         <= `ARIANE_CORE949.piton_pc_vld;
                  spc949_phy_pc_w          <= `ARIANE_CORE949.piton_pc;
                end
            end
    

            assign spc950_thread_id = 2'b00;
            assign spc950_rtl_pc = spc950_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(950*4)]   <= 1'b0;
                  active_thread[(950*4)+1] <= 1'b0;
                  active_thread[(950*4)+2] <= 1'b0;
                  active_thread[(950*4)+3] <= 1'b0;
                  spc950_inst_done         <= 0;
                  spc950_phy_pc_w          <= 0;
                end else begin
                  active_thread[(950*4)]   <= 1'b1;
                  active_thread[(950*4)+1] <= 1'b1;
                  active_thread[(950*4)+2] <= 1'b1;
                  active_thread[(950*4)+3] <= 1'b1;
                  spc950_inst_done         <= `ARIANE_CORE950.piton_pc_vld;
                  spc950_phy_pc_w          <= `ARIANE_CORE950.piton_pc;
                end
            end
    

            assign spc951_thread_id = 2'b00;
            assign spc951_rtl_pc = spc951_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(951*4)]   <= 1'b0;
                  active_thread[(951*4)+1] <= 1'b0;
                  active_thread[(951*4)+2] <= 1'b0;
                  active_thread[(951*4)+3] <= 1'b0;
                  spc951_inst_done         <= 0;
                  spc951_phy_pc_w          <= 0;
                end else begin
                  active_thread[(951*4)]   <= 1'b1;
                  active_thread[(951*4)+1] <= 1'b1;
                  active_thread[(951*4)+2] <= 1'b1;
                  active_thread[(951*4)+3] <= 1'b1;
                  spc951_inst_done         <= `ARIANE_CORE951.piton_pc_vld;
                  spc951_phy_pc_w          <= `ARIANE_CORE951.piton_pc;
                end
            end
    

            assign spc952_thread_id = 2'b00;
            assign spc952_rtl_pc = spc952_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(952*4)]   <= 1'b0;
                  active_thread[(952*4)+1] <= 1'b0;
                  active_thread[(952*4)+2] <= 1'b0;
                  active_thread[(952*4)+3] <= 1'b0;
                  spc952_inst_done         <= 0;
                  spc952_phy_pc_w          <= 0;
                end else begin
                  active_thread[(952*4)]   <= 1'b1;
                  active_thread[(952*4)+1] <= 1'b1;
                  active_thread[(952*4)+2] <= 1'b1;
                  active_thread[(952*4)+3] <= 1'b1;
                  spc952_inst_done         <= `ARIANE_CORE952.piton_pc_vld;
                  spc952_phy_pc_w          <= `ARIANE_CORE952.piton_pc;
                end
            end
    

            assign spc953_thread_id = 2'b00;
            assign spc953_rtl_pc = spc953_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(953*4)]   <= 1'b0;
                  active_thread[(953*4)+1] <= 1'b0;
                  active_thread[(953*4)+2] <= 1'b0;
                  active_thread[(953*4)+3] <= 1'b0;
                  spc953_inst_done         <= 0;
                  spc953_phy_pc_w          <= 0;
                end else begin
                  active_thread[(953*4)]   <= 1'b1;
                  active_thread[(953*4)+1] <= 1'b1;
                  active_thread[(953*4)+2] <= 1'b1;
                  active_thread[(953*4)+3] <= 1'b1;
                  spc953_inst_done         <= `ARIANE_CORE953.piton_pc_vld;
                  spc953_phy_pc_w          <= `ARIANE_CORE953.piton_pc;
                end
            end
    

            assign spc954_thread_id = 2'b00;
            assign spc954_rtl_pc = spc954_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(954*4)]   <= 1'b0;
                  active_thread[(954*4)+1] <= 1'b0;
                  active_thread[(954*4)+2] <= 1'b0;
                  active_thread[(954*4)+3] <= 1'b0;
                  spc954_inst_done         <= 0;
                  spc954_phy_pc_w          <= 0;
                end else begin
                  active_thread[(954*4)]   <= 1'b1;
                  active_thread[(954*4)+1] <= 1'b1;
                  active_thread[(954*4)+2] <= 1'b1;
                  active_thread[(954*4)+3] <= 1'b1;
                  spc954_inst_done         <= `ARIANE_CORE954.piton_pc_vld;
                  spc954_phy_pc_w          <= `ARIANE_CORE954.piton_pc;
                end
            end
    

            assign spc955_thread_id = 2'b00;
            assign spc955_rtl_pc = spc955_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(955*4)]   <= 1'b0;
                  active_thread[(955*4)+1] <= 1'b0;
                  active_thread[(955*4)+2] <= 1'b0;
                  active_thread[(955*4)+3] <= 1'b0;
                  spc955_inst_done         <= 0;
                  spc955_phy_pc_w          <= 0;
                end else begin
                  active_thread[(955*4)]   <= 1'b1;
                  active_thread[(955*4)+1] <= 1'b1;
                  active_thread[(955*4)+2] <= 1'b1;
                  active_thread[(955*4)+3] <= 1'b1;
                  spc955_inst_done         <= `ARIANE_CORE955.piton_pc_vld;
                  spc955_phy_pc_w          <= `ARIANE_CORE955.piton_pc;
                end
            end
    

            assign spc956_thread_id = 2'b00;
            assign spc956_rtl_pc = spc956_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(956*4)]   <= 1'b0;
                  active_thread[(956*4)+1] <= 1'b0;
                  active_thread[(956*4)+2] <= 1'b0;
                  active_thread[(956*4)+3] <= 1'b0;
                  spc956_inst_done         <= 0;
                  spc956_phy_pc_w          <= 0;
                end else begin
                  active_thread[(956*4)]   <= 1'b1;
                  active_thread[(956*4)+1] <= 1'b1;
                  active_thread[(956*4)+2] <= 1'b1;
                  active_thread[(956*4)+3] <= 1'b1;
                  spc956_inst_done         <= `ARIANE_CORE956.piton_pc_vld;
                  spc956_phy_pc_w          <= `ARIANE_CORE956.piton_pc;
                end
            end
    

            assign spc957_thread_id = 2'b00;
            assign spc957_rtl_pc = spc957_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(957*4)]   <= 1'b0;
                  active_thread[(957*4)+1] <= 1'b0;
                  active_thread[(957*4)+2] <= 1'b0;
                  active_thread[(957*4)+3] <= 1'b0;
                  spc957_inst_done         <= 0;
                  spc957_phy_pc_w          <= 0;
                end else begin
                  active_thread[(957*4)]   <= 1'b1;
                  active_thread[(957*4)+1] <= 1'b1;
                  active_thread[(957*4)+2] <= 1'b1;
                  active_thread[(957*4)+3] <= 1'b1;
                  spc957_inst_done         <= `ARIANE_CORE957.piton_pc_vld;
                  spc957_phy_pc_w          <= `ARIANE_CORE957.piton_pc;
                end
            end
    

            assign spc958_thread_id = 2'b00;
            assign spc958_rtl_pc = spc958_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(958*4)]   <= 1'b0;
                  active_thread[(958*4)+1] <= 1'b0;
                  active_thread[(958*4)+2] <= 1'b0;
                  active_thread[(958*4)+3] <= 1'b0;
                  spc958_inst_done         <= 0;
                  spc958_phy_pc_w          <= 0;
                end else begin
                  active_thread[(958*4)]   <= 1'b1;
                  active_thread[(958*4)+1] <= 1'b1;
                  active_thread[(958*4)+2] <= 1'b1;
                  active_thread[(958*4)+3] <= 1'b1;
                  spc958_inst_done         <= `ARIANE_CORE958.piton_pc_vld;
                  spc958_phy_pc_w          <= `ARIANE_CORE958.piton_pc;
                end
            end
    

            assign spc959_thread_id = 2'b00;
            assign spc959_rtl_pc = spc959_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(959*4)]   <= 1'b0;
                  active_thread[(959*4)+1] <= 1'b0;
                  active_thread[(959*4)+2] <= 1'b0;
                  active_thread[(959*4)+3] <= 1'b0;
                  spc959_inst_done         <= 0;
                  spc959_phy_pc_w          <= 0;
                end else begin
                  active_thread[(959*4)]   <= 1'b1;
                  active_thread[(959*4)+1] <= 1'b1;
                  active_thread[(959*4)+2] <= 1'b1;
                  active_thread[(959*4)+3] <= 1'b1;
                  spc959_inst_done         <= `ARIANE_CORE959.piton_pc_vld;
                  spc959_phy_pc_w          <= `ARIANE_CORE959.piton_pc;
                end
            end
    

            assign spc960_thread_id = 2'b00;
            assign spc960_rtl_pc = spc960_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(960*4)]   <= 1'b0;
                  active_thread[(960*4)+1] <= 1'b0;
                  active_thread[(960*4)+2] <= 1'b0;
                  active_thread[(960*4)+3] <= 1'b0;
                  spc960_inst_done         <= 0;
                  spc960_phy_pc_w          <= 0;
                end else begin
                  active_thread[(960*4)]   <= 1'b1;
                  active_thread[(960*4)+1] <= 1'b1;
                  active_thread[(960*4)+2] <= 1'b1;
                  active_thread[(960*4)+3] <= 1'b1;
                  spc960_inst_done         <= `ARIANE_CORE960.piton_pc_vld;
                  spc960_phy_pc_w          <= `ARIANE_CORE960.piton_pc;
                end
            end
    

            assign spc961_thread_id = 2'b00;
            assign spc961_rtl_pc = spc961_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(961*4)]   <= 1'b0;
                  active_thread[(961*4)+1] <= 1'b0;
                  active_thread[(961*4)+2] <= 1'b0;
                  active_thread[(961*4)+3] <= 1'b0;
                  spc961_inst_done         <= 0;
                  spc961_phy_pc_w          <= 0;
                end else begin
                  active_thread[(961*4)]   <= 1'b1;
                  active_thread[(961*4)+1] <= 1'b1;
                  active_thread[(961*4)+2] <= 1'b1;
                  active_thread[(961*4)+3] <= 1'b1;
                  spc961_inst_done         <= `ARIANE_CORE961.piton_pc_vld;
                  spc961_phy_pc_w          <= `ARIANE_CORE961.piton_pc;
                end
            end
    

            assign spc962_thread_id = 2'b00;
            assign spc962_rtl_pc = spc962_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(962*4)]   <= 1'b0;
                  active_thread[(962*4)+1] <= 1'b0;
                  active_thread[(962*4)+2] <= 1'b0;
                  active_thread[(962*4)+3] <= 1'b0;
                  spc962_inst_done         <= 0;
                  spc962_phy_pc_w          <= 0;
                end else begin
                  active_thread[(962*4)]   <= 1'b1;
                  active_thread[(962*4)+1] <= 1'b1;
                  active_thread[(962*4)+2] <= 1'b1;
                  active_thread[(962*4)+3] <= 1'b1;
                  spc962_inst_done         <= `ARIANE_CORE962.piton_pc_vld;
                  spc962_phy_pc_w          <= `ARIANE_CORE962.piton_pc;
                end
            end
    

            assign spc963_thread_id = 2'b00;
            assign spc963_rtl_pc = spc963_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(963*4)]   <= 1'b0;
                  active_thread[(963*4)+1] <= 1'b0;
                  active_thread[(963*4)+2] <= 1'b0;
                  active_thread[(963*4)+3] <= 1'b0;
                  spc963_inst_done         <= 0;
                  spc963_phy_pc_w          <= 0;
                end else begin
                  active_thread[(963*4)]   <= 1'b1;
                  active_thread[(963*4)+1] <= 1'b1;
                  active_thread[(963*4)+2] <= 1'b1;
                  active_thread[(963*4)+3] <= 1'b1;
                  spc963_inst_done         <= `ARIANE_CORE963.piton_pc_vld;
                  spc963_phy_pc_w          <= `ARIANE_CORE963.piton_pc;
                end
            end
    

            assign spc964_thread_id = 2'b00;
            assign spc964_rtl_pc = spc964_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(964*4)]   <= 1'b0;
                  active_thread[(964*4)+1] <= 1'b0;
                  active_thread[(964*4)+2] <= 1'b0;
                  active_thread[(964*4)+3] <= 1'b0;
                  spc964_inst_done         <= 0;
                  spc964_phy_pc_w          <= 0;
                end else begin
                  active_thread[(964*4)]   <= 1'b1;
                  active_thread[(964*4)+1] <= 1'b1;
                  active_thread[(964*4)+2] <= 1'b1;
                  active_thread[(964*4)+3] <= 1'b1;
                  spc964_inst_done         <= `ARIANE_CORE964.piton_pc_vld;
                  spc964_phy_pc_w          <= `ARIANE_CORE964.piton_pc;
                end
            end
    

            assign spc965_thread_id = 2'b00;
            assign spc965_rtl_pc = spc965_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(965*4)]   <= 1'b0;
                  active_thread[(965*4)+1] <= 1'b0;
                  active_thread[(965*4)+2] <= 1'b0;
                  active_thread[(965*4)+3] <= 1'b0;
                  spc965_inst_done         <= 0;
                  spc965_phy_pc_w          <= 0;
                end else begin
                  active_thread[(965*4)]   <= 1'b1;
                  active_thread[(965*4)+1] <= 1'b1;
                  active_thread[(965*4)+2] <= 1'b1;
                  active_thread[(965*4)+3] <= 1'b1;
                  spc965_inst_done         <= `ARIANE_CORE965.piton_pc_vld;
                  spc965_phy_pc_w          <= `ARIANE_CORE965.piton_pc;
                end
            end
    

            assign spc966_thread_id = 2'b00;
            assign spc966_rtl_pc = spc966_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(966*4)]   <= 1'b0;
                  active_thread[(966*4)+1] <= 1'b0;
                  active_thread[(966*4)+2] <= 1'b0;
                  active_thread[(966*4)+3] <= 1'b0;
                  spc966_inst_done         <= 0;
                  spc966_phy_pc_w          <= 0;
                end else begin
                  active_thread[(966*4)]   <= 1'b1;
                  active_thread[(966*4)+1] <= 1'b1;
                  active_thread[(966*4)+2] <= 1'b1;
                  active_thread[(966*4)+3] <= 1'b1;
                  spc966_inst_done         <= `ARIANE_CORE966.piton_pc_vld;
                  spc966_phy_pc_w          <= `ARIANE_CORE966.piton_pc;
                end
            end
    

            assign spc967_thread_id = 2'b00;
            assign spc967_rtl_pc = spc967_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(967*4)]   <= 1'b0;
                  active_thread[(967*4)+1] <= 1'b0;
                  active_thread[(967*4)+2] <= 1'b0;
                  active_thread[(967*4)+3] <= 1'b0;
                  spc967_inst_done         <= 0;
                  spc967_phy_pc_w          <= 0;
                end else begin
                  active_thread[(967*4)]   <= 1'b1;
                  active_thread[(967*4)+1] <= 1'b1;
                  active_thread[(967*4)+2] <= 1'b1;
                  active_thread[(967*4)+3] <= 1'b1;
                  spc967_inst_done         <= `ARIANE_CORE967.piton_pc_vld;
                  spc967_phy_pc_w          <= `ARIANE_CORE967.piton_pc;
                end
            end
    

            assign spc968_thread_id = 2'b00;
            assign spc968_rtl_pc = spc968_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(968*4)]   <= 1'b0;
                  active_thread[(968*4)+1] <= 1'b0;
                  active_thread[(968*4)+2] <= 1'b0;
                  active_thread[(968*4)+3] <= 1'b0;
                  spc968_inst_done         <= 0;
                  spc968_phy_pc_w          <= 0;
                end else begin
                  active_thread[(968*4)]   <= 1'b1;
                  active_thread[(968*4)+1] <= 1'b1;
                  active_thread[(968*4)+2] <= 1'b1;
                  active_thread[(968*4)+3] <= 1'b1;
                  spc968_inst_done         <= `ARIANE_CORE968.piton_pc_vld;
                  spc968_phy_pc_w          <= `ARIANE_CORE968.piton_pc;
                end
            end
    

            assign spc969_thread_id = 2'b00;
            assign spc969_rtl_pc = spc969_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(969*4)]   <= 1'b0;
                  active_thread[(969*4)+1] <= 1'b0;
                  active_thread[(969*4)+2] <= 1'b0;
                  active_thread[(969*4)+3] <= 1'b0;
                  spc969_inst_done         <= 0;
                  spc969_phy_pc_w          <= 0;
                end else begin
                  active_thread[(969*4)]   <= 1'b1;
                  active_thread[(969*4)+1] <= 1'b1;
                  active_thread[(969*4)+2] <= 1'b1;
                  active_thread[(969*4)+3] <= 1'b1;
                  spc969_inst_done         <= `ARIANE_CORE969.piton_pc_vld;
                  spc969_phy_pc_w          <= `ARIANE_CORE969.piton_pc;
                end
            end
    

            assign spc970_thread_id = 2'b00;
            assign spc970_rtl_pc = spc970_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(970*4)]   <= 1'b0;
                  active_thread[(970*4)+1] <= 1'b0;
                  active_thread[(970*4)+2] <= 1'b0;
                  active_thread[(970*4)+3] <= 1'b0;
                  spc970_inst_done         <= 0;
                  spc970_phy_pc_w          <= 0;
                end else begin
                  active_thread[(970*4)]   <= 1'b1;
                  active_thread[(970*4)+1] <= 1'b1;
                  active_thread[(970*4)+2] <= 1'b1;
                  active_thread[(970*4)+3] <= 1'b1;
                  spc970_inst_done         <= `ARIANE_CORE970.piton_pc_vld;
                  spc970_phy_pc_w          <= `ARIANE_CORE970.piton_pc;
                end
            end
    

            assign spc971_thread_id = 2'b00;
            assign spc971_rtl_pc = spc971_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(971*4)]   <= 1'b0;
                  active_thread[(971*4)+1] <= 1'b0;
                  active_thread[(971*4)+2] <= 1'b0;
                  active_thread[(971*4)+3] <= 1'b0;
                  spc971_inst_done         <= 0;
                  spc971_phy_pc_w          <= 0;
                end else begin
                  active_thread[(971*4)]   <= 1'b1;
                  active_thread[(971*4)+1] <= 1'b1;
                  active_thread[(971*4)+2] <= 1'b1;
                  active_thread[(971*4)+3] <= 1'b1;
                  spc971_inst_done         <= `ARIANE_CORE971.piton_pc_vld;
                  spc971_phy_pc_w          <= `ARIANE_CORE971.piton_pc;
                end
            end
    

            assign spc972_thread_id = 2'b00;
            assign spc972_rtl_pc = spc972_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(972*4)]   <= 1'b0;
                  active_thread[(972*4)+1] <= 1'b0;
                  active_thread[(972*4)+2] <= 1'b0;
                  active_thread[(972*4)+3] <= 1'b0;
                  spc972_inst_done         <= 0;
                  spc972_phy_pc_w          <= 0;
                end else begin
                  active_thread[(972*4)]   <= 1'b1;
                  active_thread[(972*4)+1] <= 1'b1;
                  active_thread[(972*4)+2] <= 1'b1;
                  active_thread[(972*4)+3] <= 1'b1;
                  spc972_inst_done         <= `ARIANE_CORE972.piton_pc_vld;
                  spc972_phy_pc_w          <= `ARIANE_CORE972.piton_pc;
                end
            end
    

            assign spc973_thread_id = 2'b00;
            assign spc973_rtl_pc = spc973_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(973*4)]   <= 1'b0;
                  active_thread[(973*4)+1] <= 1'b0;
                  active_thread[(973*4)+2] <= 1'b0;
                  active_thread[(973*4)+3] <= 1'b0;
                  spc973_inst_done         <= 0;
                  spc973_phy_pc_w          <= 0;
                end else begin
                  active_thread[(973*4)]   <= 1'b1;
                  active_thread[(973*4)+1] <= 1'b1;
                  active_thread[(973*4)+2] <= 1'b1;
                  active_thread[(973*4)+3] <= 1'b1;
                  spc973_inst_done         <= `ARIANE_CORE973.piton_pc_vld;
                  spc973_phy_pc_w          <= `ARIANE_CORE973.piton_pc;
                end
            end
    

            assign spc974_thread_id = 2'b00;
            assign spc974_rtl_pc = spc974_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(974*4)]   <= 1'b0;
                  active_thread[(974*4)+1] <= 1'b0;
                  active_thread[(974*4)+2] <= 1'b0;
                  active_thread[(974*4)+3] <= 1'b0;
                  spc974_inst_done         <= 0;
                  spc974_phy_pc_w          <= 0;
                end else begin
                  active_thread[(974*4)]   <= 1'b1;
                  active_thread[(974*4)+1] <= 1'b1;
                  active_thread[(974*4)+2] <= 1'b1;
                  active_thread[(974*4)+3] <= 1'b1;
                  spc974_inst_done         <= `ARIANE_CORE974.piton_pc_vld;
                  spc974_phy_pc_w          <= `ARIANE_CORE974.piton_pc;
                end
            end
    

            assign spc975_thread_id = 2'b00;
            assign spc975_rtl_pc = spc975_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(975*4)]   <= 1'b0;
                  active_thread[(975*4)+1] <= 1'b0;
                  active_thread[(975*4)+2] <= 1'b0;
                  active_thread[(975*4)+3] <= 1'b0;
                  spc975_inst_done         <= 0;
                  spc975_phy_pc_w          <= 0;
                end else begin
                  active_thread[(975*4)]   <= 1'b1;
                  active_thread[(975*4)+1] <= 1'b1;
                  active_thread[(975*4)+2] <= 1'b1;
                  active_thread[(975*4)+3] <= 1'b1;
                  spc975_inst_done         <= `ARIANE_CORE975.piton_pc_vld;
                  spc975_phy_pc_w          <= `ARIANE_CORE975.piton_pc;
                end
            end
    

            assign spc976_thread_id = 2'b00;
            assign spc976_rtl_pc = spc976_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(976*4)]   <= 1'b0;
                  active_thread[(976*4)+1] <= 1'b0;
                  active_thread[(976*4)+2] <= 1'b0;
                  active_thread[(976*4)+3] <= 1'b0;
                  spc976_inst_done         <= 0;
                  spc976_phy_pc_w          <= 0;
                end else begin
                  active_thread[(976*4)]   <= 1'b1;
                  active_thread[(976*4)+1] <= 1'b1;
                  active_thread[(976*4)+2] <= 1'b1;
                  active_thread[(976*4)+3] <= 1'b1;
                  spc976_inst_done         <= `ARIANE_CORE976.piton_pc_vld;
                  spc976_phy_pc_w          <= `ARIANE_CORE976.piton_pc;
                end
            end
    

            assign spc977_thread_id = 2'b00;
            assign spc977_rtl_pc = spc977_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(977*4)]   <= 1'b0;
                  active_thread[(977*4)+1] <= 1'b0;
                  active_thread[(977*4)+2] <= 1'b0;
                  active_thread[(977*4)+3] <= 1'b0;
                  spc977_inst_done         <= 0;
                  spc977_phy_pc_w          <= 0;
                end else begin
                  active_thread[(977*4)]   <= 1'b1;
                  active_thread[(977*4)+1] <= 1'b1;
                  active_thread[(977*4)+2] <= 1'b1;
                  active_thread[(977*4)+3] <= 1'b1;
                  spc977_inst_done         <= `ARIANE_CORE977.piton_pc_vld;
                  spc977_phy_pc_w          <= `ARIANE_CORE977.piton_pc;
                end
            end
    

            assign spc978_thread_id = 2'b00;
            assign spc978_rtl_pc = spc978_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(978*4)]   <= 1'b0;
                  active_thread[(978*4)+1] <= 1'b0;
                  active_thread[(978*4)+2] <= 1'b0;
                  active_thread[(978*4)+3] <= 1'b0;
                  spc978_inst_done         <= 0;
                  spc978_phy_pc_w          <= 0;
                end else begin
                  active_thread[(978*4)]   <= 1'b1;
                  active_thread[(978*4)+1] <= 1'b1;
                  active_thread[(978*4)+2] <= 1'b1;
                  active_thread[(978*4)+3] <= 1'b1;
                  spc978_inst_done         <= `ARIANE_CORE978.piton_pc_vld;
                  spc978_phy_pc_w          <= `ARIANE_CORE978.piton_pc;
                end
            end
    

            assign spc979_thread_id = 2'b00;
            assign spc979_rtl_pc = spc979_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(979*4)]   <= 1'b0;
                  active_thread[(979*4)+1] <= 1'b0;
                  active_thread[(979*4)+2] <= 1'b0;
                  active_thread[(979*4)+3] <= 1'b0;
                  spc979_inst_done         <= 0;
                  spc979_phy_pc_w          <= 0;
                end else begin
                  active_thread[(979*4)]   <= 1'b1;
                  active_thread[(979*4)+1] <= 1'b1;
                  active_thread[(979*4)+2] <= 1'b1;
                  active_thread[(979*4)+3] <= 1'b1;
                  spc979_inst_done         <= `ARIANE_CORE979.piton_pc_vld;
                  spc979_phy_pc_w          <= `ARIANE_CORE979.piton_pc;
                end
            end
    

            assign spc980_thread_id = 2'b00;
            assign spc980_rtl_pc = spc980_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(980*4)]   <= 1'b0;
                  active_thread[(980*4)+1] <= 1'b0;
                  active_thread[(980*4)+2] <= 1'b0;
                  active_thread[(980*4)+3] <= 1'b0;
                  spc980_inst_done         <= 0;
                  spc980_phy_pc_w          <= 0;
                end else begin
                  active_thread[(980*4)]   <= 1'b1;
                  active_thread[(980*4)+1] <= 1'b1;
                  active_thread[(980*4)+2] <= 1'b1;
                  active_thread[(980*4)+3] <= 1'b1;
                  spc980_inst_done         <= `ARIANE_CORE980.piton_pc_vld;
                  spc980_phy_pc_w          <= `ARIANE_CORE980.piton_pc;
                end
            end
    

            assign spc981_thread_id = 2'b00;
            assign spc981_rtl_pc = spc981_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(981*4)]   <= 1'b0;
                  active_thread[(981*4)+1] <= 1'b0;
                  active_thread[(981*4)+2] <= 1'b0;
                  active_thread[(981*4)+3] <= 1'b0;
                  spc981_inst_done         <= 0;
                  spc981_phy_pc_w          <= 0;
                end else begin
                  active_thread[(981*4)]   <= 1'b1;
                  active_thread[(981*4)+1] <= 1'b1;
                  active_thread[(981*4)+2] <= 1'b1;
                  active_thread[(981*4)+3] <= 1'b1;
                  spc981_inst_done         <= `ARIANE_CORE981.piton_pc_vld;
                  spc981_phy_pc_w          <= `ARIANE_CORE981.piton_pc;
                end
            end
    

            assign spc982_thread_id = 2'b00;
            assign spc982_rtl_pc = spc982_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(982*4)]   <= 1'b0;
                  active_thread[(982*4)+1] <= 1'b0;
                  active_thread[(982*4)+2] <= 1'b0;
                  active_thread[(982*4)+3] <= 1'b0;
                  spc982_inst_done         <= 0;
                  spc982_phy_pc_w          <= 0;
                end else begin
                  active_thread[(982*4)]   <= 1'b1;
                  active_thread[(982*4)+1] <= 1'b1;
                  active_thread[(982*4)+2] <= 1'b1;
                  active_thread[(982*4)+3] <= 1'b1;
                  spc982_inst_done         <= `ARIANE_CORE982.piton_pc_vld;
                  spc982_phy_pc_w          <= `ARIANE_CORE982.piton_pc;
                end
            end
    

            assign spc983_thread_id = 2'b00;
            assign spc983_rtl_pc = spc983_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(983*4)]   <= 1'b0;
                  active_thread[(983*4)+1] <= 1'b0;
                  active_thread[(983*4)+2] <= 1'b0;
                  active_thread[(983*4)+3] <= 1'b0;
                  spc983_inst_done         <= 0;
                  spc983_phy_pc_w          <= 0;
                end else begin
                  active_thread[(983*4)]   <= 1'b1;
                  active_thread[(983*4)+1] <= 1'b1;
                  active_thread[(983*4)+2] <= 1'b1;
                  active_thread[(983*4)+3] <= 1'b1;
                  spc983_inst_done         <= `ARIANE_CORE983.piton_pc_vld;
                  spc983_phy_pc_w          <= `ARIANE_CORE983.piton_pc;
                end
            end
    

            assign spc984_thread_id = 2'b00;
            assign spc984_rtl_pc = spc984_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(984*4)]   <= 1'b0;
                  active_thread[(984*4)+1] <= 1'b0;
                  active_thread[(984*4)+2] <= 1'b0;
                  active_thread[(984*4)+3] <= 1'b0;
                  spc984_inst_done         <= 0;
                  spc984_phy_pc_w          <= 0;
                end else begin
                  active_thread[(984*4)]   <= 1'b1;
                  active_thread[(984*4)+1] <= 1'b1;
                  active_thread[(984*4)+2] <= 1'b1;
                  active_thread[(984*4)+3] <= 1'b1;
                  spc984_inst_done         <= `ARIANE_CORE984.piton_pc_vld;
                  spc984_phy_pc_w          <= `ARIANE_CORE984.piton_pc;
                end
            end
    

            assign spc985_thread_id = 2'b00;
            assign spc985_rtl_pc = spc985_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(985*4)]   <= 1'b0;
                  active_thread[(985*4)+1] <= 1'b0;
                  active_thread[(985*4)+2] <= 1'b0;
                  active_thread[(985*4)+3] <= 1'b0;
                  spc985_inst_done         <= 0;
                  spc985_phy_pc_w          <= 0;
                end else begin
                  active_thread[(985*4)]   <= 1'b1;
                  active_thread[(985*4)+1] <= 1'b1;
                  active_thread[(985*4)+2] <= 1'b1;
                  active_thread[(985*4)+3] <= 1'b1;
                  spc985_inst_done         <= `ARIANE_CORE985.piton_pc_vld;
                  spc985_phy_pc_w          <= `ARIANE_CORE985.piton_pc;
                end
            end
    

            assign spc986_thread_id = 2'b00;
            assign spc986_rtl_pc = spc986_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(986*4)]   <= 1'b0;
                  active_thread[(986*4)+1] <= 1'b0;
                  active_thread[(986*4)+2] <= 1'b0;
                  active_thread[(986*4)+3] <= 1'b0;
                  spc986_inst_done         <= 0;
                  spc986_phy_pc_w          <= 0;
                end else begin
                  active_thread[(986*4)]   <= 1'b1;
                  active_thread[(986*4)+1] <= 1'b1;
                  active_thread[(986*4)+2] <= 1'b1;
                  active_thread[(986*4)+3] <= 1'b1;
                  spc986_inst_done         <= `ARIANE_CORE986.piton_pc_vld;
                  spc986_phy_pc_w          <= `ARIANE_CORE986.piton_pc;
                end
            end
    

            assign spc987_thread_id = 2'b00;
            assign spc987_rtl_pc = spc987_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(987*4)]   <= 1'b0;
                  active_thread[(987*4)+1] <= 1'b0;
                  active_thread[(987*4)+2] <= 1'b0;
                  active_thread[(987*4)+3] <= 1'b0;
                  spc987_inst_done         <= 0;
                  spc987_phy_pc_w          <= 0;
                end else begin
                  active_thread[(987*4)]   <= 1'b1;
                  active_thread[(987*4)+1] <= 1'b1;
                  active_thread[(987*4)+2] <= 1'b1;
                  active_thread[(987*4)+3] <= 1'b1;
                  spc987_inst_done         <= `ARIANE_CORE987.piton_pc_vld;
                  spc987_phy_pc_w          <= `ARIANE_CORE987.piton_pc;
                end
            end
    

            assign spc988_thread_id = 2'b00;
            assign spc988_rtl_pc = spc988_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(988*4)]   <= 1'b0;
                  active_thread[(988*4)+1] <= 1'b0;
                  active_thread[(988*4)+2] <= 1'b0;
                  active_thread[(988*4)+3] <= 1'b0;
                  spc988_inst_done         <= 0;
                  spc988_phy_pc_w          <= 0;
                end else begin
                  active_thread[(988*4)]   <= 1'b1;
                  active_thread[(988*4)+1] <= 1'b1;
                  active_thread[(988*4)+2] <= 1'b1;
                  active_thread[(988*4)+3] <= 1'b1;
                  spc988_inst_done         <= `ARIANE_CORE988.piton_pc_vld;
                  spc988_phy_pc_w          <= `ARIANE_CORE988.piton_pc;
                end
            end
    

            assign spc989_thread_id = 2'b00;
            assign spc989_rtl_pc = spc989_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(989*4)]   <= 1'b0;
                  active_thread[(989*4)+1] <= 1'b0;
                  active_thread[(989*4)+2] <= 1'b0;
                  active_thread[(989*4)+3] <= 1'b0;
                  spc989_inst_done         <= 0;
                  spc989_phy_pc_w          <= 0;
                end else begin
                  active_thread[(989*4)]   <= 1'b1;
                  active_thread[(989*4)+1] <= 1'b1;
                  active_thread[(989*4)+2] <= 1'b1;
                  active_thread[(989*4)+3] <= 1'b1;
                  spc989_inst_done         <= `ARIANE_CORE989.piton_pc_vld;
                  spc989_phy_pc_w          <= `ARIANE_CORE989.piton_pc;
                end
            end
    

            assign spc990_thread_id = 2'b00;
            assign spc990_rtl_pc = spc990_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(990*4)]   <= 1'b0;
                  active_thread[(990*4)+1] <= 1'b0;
                  active_thread[(990*4)+2] <= 1'b0;
                  active_thread[(990*4)+3] <= 1'b0;
                  spc990_inst_done         <= 0;
                  spc990_phy_pc_w          <= 0;
                end else begin
                  active_thread[(990*4)]   <= 1'b1;
                  active_thread[(990*4)+1] <= 1'b1;
                  active_thread[(990*4)+2] <= 1'b1;
                  active_thread[(990*4)+3] <= 1'b1;
                  spc990_inst_done         <= `ARIANE_CORE990.piton_pc_vld;
                  spc990_phy_pc_w          <= `ARIANE_CORE990.piton_pc;
                end
            end
    

            assign spc991_thread_id = 2'b00;
            assign spc991_rtl_pc = spc991_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(991*4)]   <= 1'b0;
                  active_thread[(991*4)+1] <= 1'b0;
                  active_thread[(991*4)+2] <= 1'b0;
                  active_thread[(991*4)+3] <= 1'b0;
                  spc991_inst_done         <= 0;
                  spc991_phy_pc_w          <= 0;
                end else begin
                  active_thread[(991*4)]   <= 1'b1;
                  active_thread[(991*4)+1] <= 1'b1;
                  active_thread[(991*4)+2] <= 1'b1;
                  active_thread[(991*4)+3] <= 1'b1;
                  spc991_inst_done         <= `ARIANE_CORE991.piton_pc_vld;
                  spc991_phy_pc_w          <= `ARIANE_CORE991.piton_pc;
                end
            end
    

            assign spc992_thread_id = 2'b00;
            assign spc992_rtl_pc = spc992_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(992*4)]   <= 1'b0;
                  active_thread[(992*4)+1] <= 1'b0;
                  active_thread[(992*4)+2] <= 1'b0;
                  active_thread[(992*4)+3] <= 1'b0;
                  spc992_inst_done         <= 0;
                  spc992_phy_pc_w          <= 0;
                end else begin
                  active_thread[(992*4)]   <= 1'b1;
                  active_thread[(992*4)+1] <= 1'b1;
                  active_thread[(992*4)+2] <= 1'b1;
                  active_thread[(992*4)+3] <= 1'b1;
                  spc992_inst_done         <= `ARIANE_CORE992.piton_pc_vld;
                  spc992_phy_pc_w          <= `ARIANE_CORE992.piton_pc;
                end
            end
    

            assign spc993_thread_id = 2'b00;
            assign spc993_rtl_pc = spc993_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(993*4)]   <= 1'b0;
                  active_thread[(993*4)+1] <= 1'b0;
                  active_thread[(993*4)+2] <= 1'b0;
                  active_thread[(993*4)+3] <= 1'b0;
                  spc993_inst_done         <= 0;
                  spc993_phy_pc_w          <= 0;
                end else begin
                  active_thread[(993*4)]   <= 1'b1;
                  active_thread[(993*4)+1] <= 1'b1;
                  active_thread[(993*4)+2] <= 1'b1;
                  active_thread[(993*4)+3] <= 1'b1;
                  spc993_inst_done         <= `ARIANE_CORE993.piton_pc_vld;
                  spc993_phy_pc_w          <= `ARIANE_CORE993.piton_pc;
                end
            end
    

            assign spc994_thread_id = 2'b00;
            assign spc994_rtl_pc = spc994_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(994*4)]   <= 1'b0;
                  active_thread[(994*4)+1] <= 1'b0;
                  active_thread[(994*4)+2] <= 1'b0;
                  active_thread[(994*4)+3] <= 1'b0;
                  spc994_inst_done         <= 0;
                  spc994_phy_pc_w          <= 0;
                end else begin
                  active_thread[(994*4)]   <= 1'b1;
                  active_thread[(994*4)+1] <= 1'b1;
                  active_thread[(994*4)+2] <= 1'b1;
                  active_thread[(994*4)+3] <= 1'b1;
                  spc994_inst_done         <= `ARIANE_CORE994.piton_pc_vld;
                  spc994_phy_pc_w          <= `ARIANE_CORE994.piton_pc;
                end
            end
    

            assign spc995_thread_id = 2'b00;
            assign spc995_rtl_pc = spc995_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(995*4)]   <= 1'b0;
                  active_thread[(995*4)+1] <= 1'b0;
                  active_thread[(995*4)+2] <= 1'b0;
                  active_thread[(995*4)+3] <= 1'b0;
                  spc995_inst_done         <= 0;
                  spc995_phy_pc_w          <= 0;
                end else begin
                  active_thread[(995*4)]   <= 1'b1;
                  active_thread[(995*4)+1] <= 1'b1;
                  active_thread[(995*4)+2] <= 1'b1;
                  active_thread[(995*4)+3] <= 1'b1;
                  spc995_inst_done         <= `ARIANE_CORE995.piton_pc_vld;
                  spc995_phy_pc_w          <= `ARIANE_CORE995.piton_pc;
                end
            end
    

            assign spc996_thread_id = 2'b00;
            assign spc996_rtl_pc = spc996_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(996*4)]   <= 1'b0;
                  active_thread[(996*4)+1] <= 1'b0;
                  active_thread[(996*4)+2] <= 1'b0;
                  active_thread[(996*4)+3] <= 1'b0;
                  spc996_inst_done         <= 0;
                  spc996_phy_pc_w          <= 0;
                end else begin
                  active_thread[(996*4)]   <= 1'b1;
                  active_thread[(996*4)+1] <= 1'b1;
                  active_thread[(996*4)+2] <= 1'b1;
                  active_thread[(996*4)+3] <= 1'b1;
                  spc996_inst_done         <= `ARIANE_CORE996.piton_pc_vld;
                  spc996_phy_pc_w          <= `ARIANE_CORE996.piton_pc;
                end
            end
    

            assign spc997_thread_id = 2'b00;
            assign spc997_rtl_pc = spc997_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(997*4)]   <= 1'b0;
                  active_thread[(997*4)+1] <= 1'b0;
                  active_thread[(997*4)+2] <= 1'b0;
                  active_thread[(997*4)+3] <= 1'b0;
                  spc997_inst_done         <= 0;
                  spc997_phy_pc_w          <= 0;
                end else begin
                  active_thread[(997*4)]   <= 1'b1;
                  active_thread[(997*4)+1] <= 1'b1;
                  active_thread[(997*4)+2] <= 1'b1;
                  active_thread[(997*4)+3] <= 1'b1;
                  spc997_inst_done         <= `ARIANE_CORE997.piton_pc_vld;
                  spc997_phy_pc_w          <= `ARIANE_CORE997.piton_pc;
                end
            end
    

            assign spc998_thread_id = 2'b00;
            assign spc998_rtl_pc = spc998_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(998*4)]   <= 1'b0;
                  active_thread[(998*4)+1] <= 1'b0;
                  active_thread[(998*4)+2] <= 1'b0;
                  active_thread[(998*4)+3] <= 1'b0;
                  spc998_inst_done         <= 0;
                  spc998_phy_pc_w          <= 0;
                end else begin
                  active_thread[(998*4)]   <= 1'b1;
                  active_thread[(998*4)+1] <= 1'b1;
                  active_thread[(998*4)+2] <= 1'b1;
                  active_thread[(998*4)+3] <= 1'b1;
                  spc998_inst_done         <= `ARIANE_CORE998.piton_pc_vld;
                  spc998_phy_pc_w          <= `ARIANE_CORE998.piton_pc;
                end
            end
    

            assign spc999_thread_id = 2'b00;
            assign spc999_rtl_pc = spc999_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(999*4)]   <= 1'b0;
                  active_thread[(999*4)+1] <= 1'b0;
                  active_thread[(999*4)+2] <= 1'b0;
                  active_thread[(999*4)+3] <= 1'b0;
                  spc999_inst_done         <= 0;
                  spc999_phy_pc_w          <= 0;
                end else begin
                  active_thread[(999*4)]   <= 1'b1;
                  active_thread[(999*4)+1] <= 1'b1;
                  active_thread[(999*4)+2] <= 1'b1;
                  active_thread[(999*4)+3] <= 1'b1;
                  spc999_inst_done         <= `ARIANE_CORE999.piton_pc_vld;
                  spc999_phy_pc_w          <= `ARIANE_CORE999.piton_pc;
                end
            end
    

            assign spc1000_thread_id = 2'b00;
            assign spc1000_rtl_pc = spc1000_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(1000*4)]   <= 1'b0;
                  active_thread[(1000*4)+1] <= 1'b0;
                  active_thread[(1000*4)+2] <= 1'b0;
                  active_thread[(1000*4)+3] <= 1'b0;
                  spc1000_inst_done         <= 0;
                  spc1000_phy_pc_w          <= 0;
                end else begin
                  active_thread[(1000*4)]   <= 1'b1;
                  active_thread[(1000*4)+1] <= 1'b1;
                  active_thread[(1000*4)+2] <= 1'b1;
                  active_thread[(1000*4)+3] <= 1'b1;
                  spc1000_inst_done         <= `ARIANE_CORE1000.piton_pc_vld;
                  spc1000_phy_pc_w          <= `ARIANE_CORE1000.piton_pc;
                end
            end
    

            assign spc1001_thread_id = 2'b00;
            assign spc1001_rtl_pc = spc1001_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(1001*4)]   <= 1'b0;
                  active_thread[(1001*4)+1] <= 1'b0;
                  active_thread[(1001*4)+2] <= 1'b0;
                  active_thread[(1001*4)+3] <= 1'b0;
                  spc1001_inst_done         <= 0;
                  spc1001_phy_pc_w          <= 0;
                end else begin
                  active_thread[(1001*4)]   <= 1'b1;
                  active_thread[(1001*4)+1] <= 1'b1;
                  active_thread[(1001*4)+2] <= 1'b1;
                  active_thread[(1001*4)+3] <= 1'b1;
                  spc1001_inst_done         <= `ARIANE_CORE1001.piton_pc_vld;
                  spc1001_phy_pc_w          <= `ARIANE_CORE1001.piton_pc;
                end
            end
    

            assign spc1002_thread_id = 2'b00;
            assign spc1002_rtl_pc = spc1002_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(1002*4)]   <= 1'b0;
                  active_thread[(1002*4)+1] <= 1'b0;
                  active_thread[(1002*4)+2] <= 1'b0;
                  active_thread[(1002*4)+3] <= 1'b0;
                  spc1002_inst_done         <= 0;
                  spc1002_phy_pc_w          <= 0;
                end else begin
                  active_thread[(1002*4)]   <= 1'b1;
                  active_thread[(1002*4)+1] <= 1'b1;
                  active_thread[(1002*4)+2] <= 1'b1;
                  active_thread[(1002*4)+3] <= 1'b1;
                  spc1002_inst_done         <= `ARIANE_CORE1002.piton_pc_vld;
                  spc1002_phy_pc_w          <= `ARIANE_CORE1002.piton_pc;
                end
            end
    

            assign spc1003_thread_id = 2'b00;
            assign spc1003_rtl_pc = spc1003_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(1003*4)]   <= 1'b0;
                  active_thread[(1003*4)+1] <= 1'b0;
                  active_thread[(1003*4)+2] <= 1'b0;
                  active_thread[(1003*4)+3] <= 1'b0;
                  spc1003_inst_done         <= 0;
                  spc1003_phy_pc_w          <= 0;
                end else begin
                  active_thread[(1003*4)]   <= 1'b1;
                  active_thread[(1003*4)+1] <= 1'b1;
                  active_thread[(1003*4)+2] <= 1'b1;
                  active_thread[(1003*4)+3] <= 1'b1;
                  spc1003_inst_done         <= `ARIANE_CORE1003.piton_pc_vld;
                  spc1003_phy_pc_w          <= `ARIANE_CORE1003.piton_pc;
                end
            end
    

            assign spc1004_thread_id = 2'b00;
            assign spc1004_rtl_pc = spc1004_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(1004*4)]   <= 1'b0;
                  active_thread[(1004*4)+1] <= 1'b0;
                  active_thread[(1004*4)+2] <= 1'b0;
                  active_thread[(1004*4)+3] <= 1'b0;
                  spc1004_inst_done         <= 0;
                  spc1004_phy_pc_w          <= 0;
                end else begin
                  active_thread[(1004*4)]   <= 1'b1;
                  active_thread[(1004*4)+1] <= 1'b1;
                  active_thread[(1004*4)+2] <= 1'b1;
                  active_thread[(1004*4)+3] <= 1'b1;
                  spc1004_inst_done         <= `ARIANE_CORE1004.piton_pc_vld;
                  spc1004_phy_pc_w          <= `ARIANE_CORE1004.piton_pc;
                end
            end
    

            assign spc1005_thread_id = 2'b00;
            assign spc1005_rtl_pc = spc1005_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(1005*4)]   <= 1'b0;
                  active_thread[(1005*4)+1] <= 1'b0;
                  active_thread[(1005*4)+2] <= 1'b0;
                  active_thread[(1005*4)+3] <= 1'b0;
                  spc1005_inst_done         <= 0;
                  spc1005_phy_pc_w          <= 0;
                end else begin
                  active_thread[(1005*4)]   <= 1'b1;
                  active_thread[(1005*4)+1] <= 1'b1;
                  active_thread[(1005*4)+2] <= 1'b1;
                  active_thread[(1005*4)+3] <= 1'b1;
                  spc1005_inst_done         <= `ARIANE_CORE1005.piton_pc_vld;
                  spc1005_phy_pc_w          <= `ARIANE_CORE1005.piton_pc;
                end
            end
    

            assign spc1006_thread_id = 2'b00;
            assign spc1006_rtl_pc = spc1006_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(1006*4)]   <= 1'b0;
                  active_thread[(1006*4)+1] <= 1'b0;
                  active_thread[(1006*4)+2] <= 1'b0;
                  active_thread[(1006*4)+3] <= 1'b0;
                  spc1006_inst_done         <= 0;
                  spc1006_phy_pc_w          <= 0;
                end else begin
                  active_thread[(1006*4)]   <= 1'b1;
                  active_thread[(1006*4)+1] <= 1'b1;
                  active_thread[(1006*4)+2] <= 1'b1;
                  active_thread[(1006*4)+3] <= 1'b1;
                  spc1006_inst_done         <= `ARIANE_CORE1006.piton_pc_vld;
                  spc1006_phy_pc_w          <= `ARIANE_CORE1006.piton_pc;
                end
            end
    

            assign spc1007_thread_id = 2'b00;
            assign spc1007_rtl_pc = spc1007_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(1007*4)]   <= 1'b0;
                  active_thread[(1007*4)+1] <= 1'b0;
                  active_thread[(1007*4)+2] <= 1'b0;
                  active_thread[(1007*4)+3] <= 1'b0;
                  spc1007_inst_done         <= 0;
                  spc1007_phy_pc_w          <= 0;
                end else begin
                  active_thread[(1007*4)]   <= 1'b1;
                  active_thread[(1007*4)+1] <= 1'b1;
                  active_thread[(1007*4)+2] <= 1'b1;
                  active_thread[(1007*4)+3] <= 1'b1;
                  spc1007_inst_done         <= `ARIANE_CORE1007.piton_pc_vld;
                  spc1007_phy_pc_w          <= `ARIANE_CORE1007.piton_pc;
                end
            end
    

            assign spc1008_thread_id = 2'b00;
            assign spc1008_rtl_pc = spc1008_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(1008*4)]   <= 1'b0;
                  active_thread[(1008*4)+1] <= 1'b0;
                  active_thread[(1008*4)+2] <= 1'b0;
                  active_thread[(1008*4)+3] <= 1'b0;
                  spc1008_inst_done         <= 0;
                  spc1008_phy_pc_w          <= 0;
                end else begin
                  active_thread[(1008*4)]   <= 1'b1;
                  active_thread[(1008*4)+1] <= 1'b1;
                  active_thread[(1008*4)+2] <= 1'b1;
                  active_thread[(1008*4)+3] <= 1'b1;
                  spc1008_inst_done         <= `ARIANE_CORE1008.piton_pc_vld;
                  spc1008_phy_pc_w          <= `ARIANE_CORE1008.piton_pc;
                end
            end
    

            assign spc1009_thread_id = 2'b00;
            assign spc1009_rtl_pc = spc1009_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(1009*4)]   <= 1'b0;
                  active_thread[(1009*4)+1] <= 1'b0;
                  active_thread[(1009*4)+2] <= 1'b0;
                  active_thread[(1009*4)+3] <= 1'b0;
                  spc1009_inst_done         <= 0;
                  spc1009_phy_pc_w          <= 0;
                end else begin
                  active_thread[(1009*4)]   <= 1'b1;
                  active_thread[(1009*4)+1] <= 1'b1;
                  active_thread[(1009*4)+2] <= 1'b1;
                  active_thread[(1009*4)+3] <= 1'b1;
                  spc1009_inst_done         <= `ARIANE_CORE1009.piton_pc_vld;
                  spc1009_phy_pc_w          <= `ARIANE_CORE1009.piton_pc;
                end
            end
    

            assign spc1010_thread_id = 2'b00;
            assign spc1010_rtl_pc = spc1010_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(1010*4)]   <= 1'b0;
                  active_thread[(1010*4)+1] <= 1'b0;
                  active_thread[(1010*4)+2] <= 1'b0;
                  active_thread[(1010*4)+3] <= 1'b0;
                  spc1010_inst_done         <= 0;
                  spc1010_phy_pc_w          <= 0;
                end else begin
                  active_thread[(1010*4)]   <= 1'b1;
                  active_thread[(1010*4)+1] <= 1'b1;
                  active_thread[(1010*4)+2] <= 1'b1;
                  active_thread[(1010*4)+3] <= 1'b1;
                  spc1010_inst_done         <= `ARIANE_CORE1010.piton_pc_vld;
                  spc1010_phy_pc_w          <= `ARIANE_CORE1010.piton_pc;
                end
            end
    

            assign spc1011_thread_id = 2'b00;
            assign spc1011_rtl_pc = spc1011_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(1011*4)]   <= 1'b0;
                  active_thread[(1011*4)+1] <= 1'b0;
                  active_thread[(1011*4)+2] <= 1'b0;
                  active_thread[(1011*4)+3] <= 1'b0;
                  spc1011_inst_done         <= 0;
                  spc1011_phy_pc_w          <= 0;
                end else begin
                  active_thread[(1011*4)]   <= 1'b1;
                  active_thread[(1011*4)+1] <= 1'b1;
                  active_thread[(1011*4)+2] <= 1'b1;
                  active_thread[(1011*4)+3] <= 1'b1;
                  spc1011_inst_done         <= `ARIANE_CORE1011.piton_pc_vld;
                  spc1011_phy_pc_w          <= `ARIANE_CORE1011.piton_pc;
                end
            end
    

            assign spc1012_thread_id = 2'b00;
            assign spc1012_rtl_pc = spc1012_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(1012*4)]   <= 1'b0;
                  active_thread[(1012*4)+1] <= 1'b0;
                  active_thread[(1012*4)+2] <= 1'b0;
                  active_thread[(1012*4)+3] <= 1'b0;
                  spc1012_inst_done         <= 0;
                  spc1012_phy_pc_w          <= 0;
                end else begin
                  active_thread[(1012*4)]   <= 1'b1;
                  active_thread[(1012*4)+1] <= 1'b1;
                  active_thread[(1012*4)+2] <= 1'b1;
                  active_thread[(1012*4)+3] <= 1'b1;
                  spc1012_inst_done         <= `ARIANE_CORE1012.piton_pc_vld;
                  spc1012_phy_pc_w          <= `ARIANE_CORE1012.piton_pc;
                end
            end
    

            assign spc1013_thread_id = 2'b00;
            assign spc1013_rtl_pc = spc1013_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(1013*4)]   <= 1'b0;
                  active_thread[(1013*4)+1] <= 1'b0;
                  active_thread[(1013*4)+2] <= 1'b0;
                  active_thread[(1013*4)+3] <= 1'b0;
                  spc1013_inst_done         <= 0;
                  spc1013_phy_pc_w          <= 0;
                end else begin
                  active_thread[(1013*4)]   <= 1'b1;
                  active_thread[(1013*4)+1] <= 1'b1;
                  active_thread[(1013*4)+2] <= 1'b1;
                  active_thread[(1013*4)+3] <= 1'b1;
                  spc1013_inst_done         <= `ARIANE_CORE1013.piton_pc_vld;
                  spc1013_phy_pc_w          <= `ARIANE_CORE1013.piton_pc;
                end
            end
    

            assign spc1014_thread_id = 2'b00;
            assign spc1014_rtl_pc = spc1014_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(1014*4)]   <= 1'b0;
                  active_thread[(1014*4)+1] <= 1'b0;
                  active_thread[(1014*4)+2] <= 1'b0;
                  active_thread[(1014*4)+3] <= 1'b0;
                  spc1014_inst_done         <= 0;
                  spc1014_phy_pc_w          <= 0;
                end else begin
                  active_thread[(1014*4)]   <= 1'b1;
                  active_thread[(1014*4)+1] <= 1'b1;
                  active_thread[(1014*4)+2] <= 1'b1;
                  active_thread[(1014*4)+3] <= 1'b1;
                  spc1014_inst_done         <= `ARIANE_CORE1014.piton_pc_vld;
                  spc1014_phy_pc_w          <= `ARIANE_CORE1014.piton_pc;
                end
            end
    

            assign spc1015_thread_id = 2'b00;
            assign spc1015_rtl_pc = spc1015_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(1015*4)]   <= 1'b0;
                  active_thread[(1015*4)+1] <= 1'b0;
                  active_thread[(1015*4)+2] <= 1'b0;
                  active_thread[(1015*4)+3] <= 1'b0;
                  spc1015_inst_done         <= 0;
                  spc1015_phy_pc_w          <= 0;
                end else begin
                  active_thread[(1015*4)]   <= 1'b1;
                  active_thread[(1015*4)+1] <= 1'b1;
                  active_thread[(1015*4)+2] <= 1'b1;
                  active_thread[(1015*4)+3] <= 1'b1;
                  spc1015_inst_done         <= `ARIANE_CORE1015.piton_pc_vld;
                  spc1015_phy_pc_w          <= `ARIANE_CORE1015.piton_pc;
                end
            end
    

            assign spc1016_thread_id = 2'b00;
            assign spc1016_rtl_pc = spc1016_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(1016*4)]   <= 1'b0;
                  active_thread[(1016*4)+1] <= 1'b0;
                  active_thread[(1016*4)+2] <= 1'b0;
                  active_thread[(1016*4)+3] <= 1'b0;
                  spc1016_inst_done         <= 0;
                  spc1016_phy_pc_w          <= 0;
                end else begin
                  active_thread[(1016*4)]   <= 1'b1;
                  active_thread[(1016*4)+1] <= 1'b1;
                  active_thread[(1016*4)+2] <= 1'b1;
                  active_thread[(1016*4)+3] <= 1'b1;
                  spc1016_inst_done         <= `ARIANE_CORE1016.piton_pc_vld;
                  spc1016_phy_pc_w          <= `ARIANE_CORE1016.piton_pc;
                end
            end
    

            assign spc1017_thread_id = 2'b00;
            assign spc1017_rtl_pc = spc1017_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(1017*4)]   <= 1'b0;
                  active_thread[(1017*4)+1] <= 1'b0;
                  active_thread[(1017*4)+2] <= 1'b0;
                  active_thread[(1017*4)+3] <= 1'b0;
                  spc1017_inst_done         <= 0;
                  spc1017_phy_pc_w          <= 0;
                end else begin
                  active_thread[(1017*4)]   <= 1'b1;
                  active_thread[(1017*4)+1] <= 1'b1;
                  active_thread[(1017*4)+2] <= 1'b1;
                  active_thread[(1017*4)+3] <= 1'b1;
                  spc1017_inst_done         <= `ARIANE_CORE1017.piton_pc_vld;
                  spc1017_phy_pc_w          <= `ARIANE_CORE1017.piton_pc;
                end
            end
    

            assign spc1018_thread_id = 2'b00;
            assign spc1018_rtl_pc = spc1018_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(1018*4)]   <= 1'b0;
                  active_thread[(1018*4)+1] <= 1'b0;
                  active_thread[(1018*4)+2] <= 1'b0;
                  active_thread[(1018*4)+3] <= 1'b0;
                  spc1018_inst_done         <= 0;
                  spc1018_phy_pc_w          <= 0;
                end else begin
                  active_thread[(1018*4)]   <= 1'b1;
                  active_thread[(1018*4)+1] <= 1'b1;
                  active_thread[(1018*4)+2] <= 1'b1;
                  active_thread[(1018*4)+3] <= 1'b1;
                  spc1018_inst_done         <= `ARIANE_CORE1018.piton_pc_vld;
                  spc1018_phy_pc_w          <= `ARIANE_CORE1018.piton_pc;
                end
            end
    

            assign spc1019_thread_id = 2'b00;
            assign spc1019_rtl_pc = spc1019_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(1019*4)]   <= 1'b0;
                  active_thread[(1019*4)+1] <= 1'b0;
                  active_thread[(1019*4)+2] <= 1'b0;
                  active_thread[(1019*4)+3] <= 1'b0;
                  spc1019_inst_done         <= 0;
                  spc1019_phy_pc_w          <= 0;
                end else begin
                  active_thread[(1019*4)]   <= 1'b1;
                  active_thread[(1019*4)+1] <= 1'b1;
                  active_thread[(1019*4)+2] <= 1'b1;
                  active_thread[(1019*4)+3] <= 1'b1;
                  spc1019_inst_done         <= `ARIANE_CORE1019.piton_pc_vld;
                  spc1019_phy_pc_w          <= `ARIANE_CORE1019.piton_pc;
                end
            end
    

            assign spc1020_thread_id = 2'b00;
            assign spc1020_rtl_pc = spc1020_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(1020*4)]   <= 1'b0;
                  active_thread[(1020*4)+1] <= 1'b0;
                  active_thread[(1020*4)+2] <= 1'b0;
                  active_thread[(1020*4)+3] <= 1'b0;
                  spc1020_inst_done         <= 0;
                  spc1020_phy_pc_w          <= 0;
                end else begin
                  active_thread[(1020*4)]   <= 1'b1;
                  active_thread[(1020*4)+1] <= 1'b1;
                  active_thread[(1020*4)+2] <= 1'b1;
                  active_thread[(1020*4)+3] <= 1'b1;
                  spc1020_inst_done         <= `ARIANE_CORE1020.piton_pc_vld;
                  spc1020_phy_pc_w          <= `ARIANE_CORE1020.piton_pc;
                end
            end
    

            assign spc1021_thread_id = 2'b00;
            assign spc1021_rtl_pc = spc1021_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(1021*4)]   <= 1'b0;
                  active_thread[(1021*4)+1] <= 1'b0;
                  active_thread[(1021*4)+2] <= 1'b0;
                  active_thread[(1021*4)+3] <= 1'b0;
                  spc1021_inst_done         <= 0;
                  spc1021_phy_pc_w          <= 0;
                end else begin
                  active_thread[(1021*4)]   <= 1'b1;
                  active_thread[(1021*4)+1] <= 1'b1;
                  active_thread[(1021*4)+2] <= 1'b1;
                  active_thread[(1021*4)+3] <= 1'b1;
                  spc1021_inst_done         <= `ARIANE_CORE1021.piton_pc_vld;
                  spc1021_phy_pc_w          <= `ARIANE_CORE1021.piton_pc;
                end
            end
    

            assign spc1022_thread_id = 2'b00;
            assign spc1022_rtl_pc = spc1022_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(1022*4)]   <= 1'b0;
                  active_thread[(1022*4)+1] <= 1'b0;
                  active_thread[(1022*4)+2] <= 1'b0;
                  active_thread[(1022*4)+3] <= 1'b0;
                  spc1022_inst_done         <= 0;
                  spc1022_phy_pc_w          <= 0;
                end else begin
                  active_thread[(1022*4)]   <= 1'b1;
                  active_thread[(1022*4)+1] <= 1'b1;
                  active_thread[(1022*4)+2] <= 1'b1;
                  active_thread[(1022*4)+3] <= 1'b1;
                  spc1022_inst_done         <= `ARIANE_CORE1022.piton_pc_vld;
                  spc1022_phy_pc_w          <= `ARIANE_CORE1022.piton_pc;
                end
            end
    

            assign spc1023_thread_id = 2'b00;
            assign spc1023_rtl_pc = spc1023_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(1023*4)]   <= 1'b0;
                  active_thread[(1023*4)+1] <= 1'b0;
                  active_thread[(1023*4)+2] <= 1'b0;
                  active_thread[(1023*4)+3] <= 1'b0;
                  spc1023_inst_done         <= 0;
                  spc1023_phy_pc_w          <= 0;
                end else begin
                  active_thread[(1023*4)]   <= 1'b1;
                  active_thread[(1023*4)+1] <= 1'b1;
                  active_thread[(1023*4)+2] <= 1'b1;
                  active_thread[(1023*4)+3] <= 1'b1;
                  spc1023_inst_done         <= `ARIANE_CORE1023.piton_pc_vld;
                  spc1023_phy_pc_w          <= `ARIANE_CORE1023.piton_pc;
                end
            end
    




reg           dummy;

task trap_extract;
    reg [2048:0] pc_str;
    reg [63:0]  tmp_val;
    integer     i;
    begin
        bad_trap_count = 0;

            if($value$plusargs("good_trap0=%h", tmp_val)) begin
                good_trap[0] = tmp_val;
                good_trap_exists[0] = 1'b1;
                //$display ("%t: good_trap %h", $time, good_trap[0]);
            end



            if($value$plusargs("bad_trap0=%h", tmp_val)) begin
                bad_trap[0] = tmp_val;
                bad_trap_exists[0] = 1'b1;
                //$display ("%t: bad_trap %h", $time, bad_trap[0]);
            end

        trap_count = good_trap_count > bad_trap_count ? good_trap_count :  bad_trap_count;

    end
endtask // trap_extract
// deceide pass or fail
integer       ind;
//post-silicon request
reg [63:0]    last_hit [31:0];
//indicate the 2nd time hit.
reg [31:0]    hitted;
initial hitted = 0;

reg first_rst;
initial begin
    //#20//need to wait for socket initializing.
     trap_extract;
    done    = 0;
    first_rst = 1;
    for(ind = 0;ind < `PITON_NUM_TILES; ind = ind + 1)timeout[ind] = 0;
end // initial begin
always @(posedge rst_l)begin
    if(first_rst)begin
        active_thread = 0;
        first_rst     = 0;
        done          = 0;
    end
end

task set_diag_done;
    input local_diag_done;

    begin
        if (local_diag_done) begin
            `TOP_MOD.diag_done = 1;
        end
    end
endtask


    wire[31:0] long_cpuid0;
    assign long_cpuid0 = {30'd0, spc0_thread_id};

    wire[31:0] long_cpuid1;
    assign long_cpuid1 = {30'd1, spc1_thread_id};

    wire[31:0] long_cpuid2;
    assign long_cpuid2 = {30'd2, spc2_thread_id};

    wire[31:0] long_cpuid3;
    assign long_cpuid3 = {30'd3, spc3_thread_id};

    wire[31:0] long_cpuid4;
    assign long_cpuid4 = {30'd4, spc4_thread_id};

    wire[31:0] long_cpuid5;
    assign long_cpuid5 = {30'd5, spc5_thread_id};

    wire[31:0] long_cpuid6;
    assign long_cpuid6 = {30'd6, spc6_thread_id};

    wire[31:0] long_cpuid7;
    assign long_cpuid7 = {30'd7, spc7_thread_id};

    wire[31:0] long_cpuid8;
    assign long_cpuid8 = {30'd8, spc8_thread_id};

    wire[31:0] long_cpuid9;
    assign long_cpuid9 = {30'd9, spc9_thread_id};

    wire[31:0] long_cpuid10;
    assign long_cpuid10 = {30'd10, spc10_thread_id};

    wire[31:0] long_cpuid11;
    assign long_cpuid11 = {30'd11, spc11_thread_id};

    wire[31:0] long_cpuid12;
    assign long_cpuid12 = {30'd12, spc12_thread_id};

    wire[31:0] long_cpuid13;
    assign long_cpuid13 = {30'd13, spc13_thread_id};

    wire[31:0] long_cpuid14;
    assign long_cpuid14 = {30'd14, spc14_thread_id};

    wire[31:0] long_cpuid15;
    assign long_cpuid15 = {30'd15, spc15_thread_id};

    wire[31:0] long_cpuid16;
    assign long_cpuid16 = {30'd16, spc16_thread_id};

    wire[31:0] long_cpuid17;
    assign long_cpuid17 = {30'd17, spc17_thread_id};

    wire[31:0] long_cpuid18;
    assign long_cpuid18 = {30'd18, spc18_thread_id};

    wire[31:0] long_cpuid19;
    assign long_cpuid19 = {30'd19, spc19_thread_id};

    wire[31:0] long_cpuid20;
    assign long_cpuid20 = {30'd20, spc20_thread_id};

    wire[31:0] long_cpuid21;
    assign long_cpuid21 = {30'd21, spc21_thread_id};

    wire[31:0] long_cpuid22;
    assign long_cpuid22 = {30'd22, spc22_thread_id};

    wire[31:0] long_cpuid23;
    assign long_cpuid23 = {30'd23, spc23_thread_id};

    wire[31:0] long_cpuid24;
    assign long_cpuid24 = {30'd24, spc24_thread_id};

    wire[31:0] long_cpuid25;
    assign long_cpuid25 = {30'd25, spc25_thread_id};

    wire[31:0] long_cpuid26;
    assign long_cpuid26 = {30'd26, spc26_thread_id};

    wire[31:0] long_cpuid27;
    assign long_cpuid27 = {30'd27, spc27_thread_id};

    wire[31:0] long_cpuid28;
    assign long_cpuid28 = {30'd28, spc28_thread_id};

    wire[31:0] long_cpuid29;
    assign long_cpuid29 = {30'd29, spc29_thread_id};

    wire[31:0] long_cpuid30;
    assign long_cpuid30 = {30'd30, spc30_thread_id};

    wire[31:0] long_cpuid31;
    assign long_cpuid31 = {30'd31, spc31_thread_id};

    wire[31:0] long_cpuid32;
    assign long_cpuid32 = {30'd32, spc32_thread_id};

    wire[31:0] long_cpuid33;
    assign long_cpuid33 = {30'd33, spc33_thread_id};

    wire[31:0] long_cpuid34;
    assign long_cpuid34 = {30'd34, spc34_thread_id};

    wire[31:0] long_cpuid35;
    assign long_cpuid35 = {30'd35, spc35_thread_id};

    wire[31:0] long_cpuid36;
    assign long_cpuid36 = {30'd36, spc36_thread_id};

    wire[31:0] long_cpuid37;
    assign long_cpuid37 = {30'd37, spc37_thread_id};

    wire[31:0] long_cpuid38;
    assign long_cpuid38 = {30'd38, spc38_thread_id};

    wire[31:0] long_cpuid39;
    assign long_cpuid39 = {30'd39, spc39_thread_id};

    wire[31:0] long_cpuid40;
    assign long_cpuid40 = {30'd40, spc40_thread_id};

    wire[31:0] long_cpuid41;
    assign long_cpuid41 = {30'd41, spc41_thread_id};

    wire[31:0] long_cpuid42;
    assign long_cpuid42 = {30'd42, spc42_thread_id};

    wire[31:0] long_cpuid43;
    assign long_cpuid43 = {30'd43, spc43_thread_id};

    wire[31:0] long_cpuid44;
    assign long_cpuid44 = {30'd44, spc44_thread_id};

    wire[31:0] long_cpuid45;
    assign long_cpuid45 = {30'd45, spc45_thread_id};

    wire[31:0] long_cpuid46;
    assign long_cpuid46 = {30'd46, spc46_thread_id};

    wire[31:0] long_cpuid47;
    assign long_cpuid47 = {30'd47, spc47_thread_id};

    wire[31:0] long_cpuid48;
    assign long_cpuid48 = {30'd48, spc48_thread_id};

    wire[31:0] long_cpuid49;
    assign long_cpuid49 = {30'd49, spc49_thread_id};

    wire[31:0] long_cpuid50;
    assign long_cpuid50 = {30'd50, spc50_thread_id};

    wire[31:0] long_cpuid51;
    assign long_cpuid51 = {30'd51, spc51_thread_id};

    wire[31:0] long_cpuid52;
    assign long_cpuid52 = {30'd52, spc52_thread_id};

    wire[31:0] long_cpuid53;
    assign long_cpuid53 = {30'd53, spc53_thread_id};

    wire[31:0] long_cpuid54;
    assign long_cpuid54 = {30'd54, spc54_thread_id};

    wire[31:0] long_cpuid55;
    assign long_cpuid55 = {30'd55, spc55_thread_id};

    wire[31:0] long_cpuid56;
    assign long_cpuid56 = {30'd56, spc56_thread_id};

    wire[31:0] long_cpuid57;
    assign long_cpuid57 = {30'd57, spc57_thread_id};

    wire[31:0] long_cpuid58;
    assign long_cpuid58 = {30'd58, spc58_thread_id};

    wire[31:0] long_cpuid59;
    assign long_cpuid59 = {30'd59, spc59_thread_id};

    wire[31:0] long_cpuid60;
    assign long_cpuid60 = {30'd60, spc60_thread_id};

    wire[31:0] long_cpuid61;
    assign long_cpuid61 = {30'd61, spc61_thread_id};

    wire[31:0] long_cpuid62;
    assign long_cpuid62 = {30'd62, spc62_thread_id};

    wire[31:0] long_cpuid63;
    assign long_cpuid63 = {30'd63, spc63_thread_id};

    wire[31:0] long_cpuid64;
    assign long_cpuid64 = {30'd64, spc64_thread_id};

    wire[31:0] long_cpuid65;
    assign long_cpuid65 = {30'd65, spc65_thread_id};

    wire[31:0] long_cpuid66;
    assign long_cpuid66 = {30'd66, spc66_thread_id};

    wire[31:0] long_cpuid67;
    assign long_cpuid67 = {30'd67, spc67_thread_id};

    wire[31:0] long_cpuid68;
    assign long_cpuid68 = {30'd68, spc68_thread_id};

    wire[31:0] long_cpuid69;
    assign long_cpuid69 = {30'd69, spc69_thread_id};

    wire[31:0] long_cpuid70;
    assign long_cpuid70 = {30'd70, spc70_thread_id};

    wire[31:0] long_cpuid71;
    assign long_cpuid71 = {30'd71, spc71_thread_id};

    wire[31:0] long_cpuid72;
    assign long_cpuid72 = {30'd72, spc72_thread_id};

    wire[31:0] long_cpuid73;
    assign long_cpuid73 = {30'd73, spc73_thread_id};

    wire[31:0] long_cpuid74;
    assign long_cpuid74 = {30'd74, spc74_thread_id};

    wire[31:0] long_cpuid75;
    assign long_cpuid75 = {30'd75, spc75_thread_id};

    wire[31:0] long_cpuid76;
    assign long_cpuid76 = {30'd76, spc76_thread_id};

    wire[31:0] long_cpuid77;
    assign long_cpuid77 = {30'd77, spc77_thread_id};

    wire[31:0] long_cpuid78;
    assign long_cpuid78 = {30'd78, spc78_thread_id};

    wire[31:0] long_cpuid79;
    assign long_cpuid79 = {30'd79, spc79_thread_id};

    wire[31:0] long_cpuid80;
    assign long_cpuid80 = {30'd80, spc80_thread_id};

    wire[31:0] long_cpuid81;
    assign long_cpuid81 = {30'd81, spc81_thread_id};

    wire[31:0] long_cpuid82;
    assign long_cpuid82 = {30'd82, spc82_thread_id};

    wire[31:0] long_cpuid83;
    assign long_cpuid83 = {30'd83, spc83_thread_id};

    wire[31:0] long_cpuid84;
    assign long_cpuid84 = {30'd84, spc84_thread_id};

    wire[31:0] long_cpuid85;
    assign long_cpuid85 = {30'd85, spc85_thread_id};

    wire[31:0] long_cpuid86;
    assign long_cpuid86 = {30'd86, spc86_thread_id};

    wire[31:0] long_cpuid87;
    assign long_cpuid87 = {30'd87, spc87_thread_id};

    wire[31:0] long_cpuid88;
    assign long_cpuid88 = {30'd88, spc88_thread_id};

    wire[31:0] long_cpuid89;
    assign long_cpuid89 = {30'd89, spc89_thread_id};

    wire[31:0] long_cpuid90;
    assign long_cpuid90 = {30'd90, spc90_thread_id};

    wire[31:0] long_cpuid91;
    assign long_cpuid91 = {30'd91, spc91_thread_id};

    wire[31:0] long_cpuid92;
    assign long_cpuid92 = {30'd92, spc92_thread_id};

    wire[31:0] long_cpuid93;
    assign long_cpuid93 = {30'd93, spc93_thread_id};

    wire[31:0] long_cpuid94;
    assign long_cpuid94 = {30'd94, spc94_thread_id};

    wire[31:0] long_cpuid95;
    assign long_cpuid95 = {30'd95, spc95_thread_id};

    wire[31:0] long_cpuid96;
    assign long_cpuid96 = {30'd96, spc96_thread_id};

    wire[31:0] long_cpuid97;
    assign long_cpuid97 = {30'd97, spc97_thread_id};

    wire[31:0] long_cpuid98;
    assign long_cpuid98 = {30'd98, spc98_thread_id};

    wire[31:0] long_cpuid99;
    assign long_cpuid99 = {30'd99, spc99_thread_id};

    wire[31:0] long_cpuid100;
    assign long_cpuid100 = {30'd100, spc100_thread_id};

    wire[31:0] long_cpuid101;
    assign long_cpuid101 = {30'd101, spc101_thread_id};

    wire[31:0] long_cpuid102;
    assign long_cpuid102 = {30'd102, spc102_thread_id};

    wire[31:0] long_cpuid103;
    assign long_cpuid103 = {30'd103, spc103_thread_id};

    wire[31:0] long_cpuid104;
    assign long_cpuid104 = {30'd104, spc104_thread_id};

    wire[31:0] long_cpuid105;
    assign long_cpuid105 = {30'd105, spc105_thread_id};

    wire[31:0] long_cpuid106;
    assign long_cpuid106 = {30'd106, spc106_thread_id};

    wire[31:0] long_cpuid107;
    assign long_cpuid107 = {30'd107, spc107_thread_id};

    wire[31:0] long_cpuid108;
    assign long_cpuid108 = {30'd108, spc108_thread_id};

    wire[31:0] long_cpuid109;
    assign long_cpuid109 = {30'd109, spc109_thread_id};

    wire[31:0] long_cpuid110;
    assign long_cpuid110 = {30'd110, spc110_thread_id};

    wire[31:0] long_cpuid111;
    assign long_cpuid111 = {30'd111, spc111_thread_id};

    wire[31:0] long_cpuid112;
    assign long_cpuid112 = {30'd112, spc112_thread_id};

    wire[31:0] long_cpuid113;
    assign long_cpuid113 = {30'd113, spc113_thread_id};

    wire[31:0] long_cpuid114;
    assign long_cpuid114 = {30'd114, spc114_thread_id};

    wire[31:0] long_cpuid115;
    assign long_cpuid115 = {30'd115, spc115_thread_id};

    wire[31:0] long_cpuid116;
    assign long_cpuid116 = {30'd116, spc116_thread_id};

    wire[31:0] long_cpuid117;
    assign long_cpuid117 = {30'd117, spc117_thread_id};

    wire[31:0] long_cpuid118;
    assign long_cpuid118 = {30'd118, spc118_thread_id};

    wire[31:0] long_cpuid119;
    assign long_cpuid119 = {30'd119, spc119_thread_id};

    wire[31:0] long_cpuid120;
    assign long_cpuid120 = {30'd120, spc120_thread_id};

    wire[31:0] long_cpuid121;
    assign long_cpuid121 = {30'd121, spc121_thread_id};

    wire[31:0] long_cpuid122;
    assign long_cpuid122 = {30'd122, spc122_thread_id};

    wire[31:0] long_cpuid123;
    assign long_cpuid123 = {30'd123, spc123_thread_id};

    wire[31:0] long_cpuid124;
    assign long_cpuid124 = {30'd124, spc124_thread_id};

    wire[31:0] long_cpuid125;
    assign long_cpuid125 = {30'd125, spc125_thread_id};

    wire[31:0] long_cpuid126;
    assign long_cpuid126 = {30'd126, spc126_thread_id};

    wire[31:0] long_cpuid127;
    assign long_cpuid127 = {30'd127, spc127_thread_id};

    wire[31:0] long_cpuid128;
    assign long_cpuid128 = {30'd128, spc128_thread_id};

    wire[31:0] long_cpuid129;
    assign long_cpuid129 = {30'd129, spc129_thread_id};

    wire[31:0] long_cpuid130;
    assign long_cpuid130 = {30'd130, spc130_thread_id};

    wire[31:0] long_cpuid131;
    assign long_cpuid131 = {30'd131, spc131_thread_id};

    wire[31:0] long_cpuid132;
    assign long_cpuid132 = {30'd132, spc132_thread_id};

    wire[31:0] long_cpuid133;
    assign long_cpuid133 = {30'd133, spc133_thread_id};

    wire[31:0] long_cpuid134;
    assign long_cpuid134 = {30'd134, spc134_thread_id};

    wire[31:0] long_cpuid135;
    assign long_cpuid135 = {30'd135, spc135_thread_id};

    wire[31:0] long_cpuid136;
    assign long_cpuid136 = {30'd136, spc136_thread_id};

    wire[31:0] long_cpuid137;
    assign long_cpuid137 = {30'd137, spc137_thread_id};

    wire[31:0] long_cpuid138;
    assign long_cpuid138 = {30'd138, spc138_thread_id};

    wire[31:0] long_cpuid139;
    assign long_cpuid139 = {30'd139, spc139_thread_id};

    wire[31:0] long_cpuid140;
    assign long_cpuid140 = {30'd140, spc140_thread_id};

    wire[31:0] long_cpuid141;
    assign long_cpuid141 = {30'd141, spc141_thread_id};

    wire[31:0] long_cpuid142;
    assign long_cpuid142 = {30'd142, spc142_thread_id};

    wire[31:0] long_cpuid143;
    assign long_cpuid143 = {30'd143, spc143_thread_id};

    wire[31:0] long_cpuid144;
    assign long_cpuid144 = {30'd144, spc144_thread_id};

    wire[31:0] long_cpuid145;
    assign long_cpuid145 = {30'd145, spc145_thread_id};

    wire[31:0] long_cpuid146;
    assign long_cpuid146 = {30'd146, spc146_thread_id};

    wire[31:0] long_cpuid147;
    assign long_cpuid147 = {30'd147, spc147_thread_id};

    wire[31:0] long_cpuid148;
    assign long_cpuid148 = {30'd148, spc148_thread_id};

    wire[31:0] long_cpuid149;
    assign long_cpuid149 = {30'd149, spc149_thread_id};

    wire[31:0] long_cpuid150;
    assign long_cpuid150 = {30'd150, spc150_thread_id};

    wire[31:0] long_cpuid151;
    assign long_cpuid151 = {30'd151, spc151_thread_id};

    wire[31:0] long_cpuid152;
    assign long_cpuid152 = {30'd152, spc152_thread_id};

    wire[31:0] long_cpuid153;
    assign long_cpuid153 = {30'd153, spc153_thread_id};

    wire[31:0] long_cpuid154;
    assign long_cpuid154 = {30'd154, spc154_thread_id};

    wire[31:0] long_cpuid155;
    assign long_cpuid155 = {30'd155, spc155_thread_id};

    wire[31:0] long_cpuid156;
    assign long_cpuid156 = {30'd156, spc156_thread_id};

    wire[31:0] long_cpuid157;
    assign long_cpuid157 = {30'd157, spc157_thread_id};

    wire[31:0] long_cpuid158;
    assign long_cpuid158 = {30'd158, spc158_thread_id};

    wire[31:0] long_cpuid159;
    assign long_cpuid159 = {30'd159, spc159_thread_id};

    wire[31:0] long_cpuid160;
    assign long_cpuid160 = {30'd160, spc160_thread_id};

    wire[31:0] long_cpuid161;
    assign long_cpuid161 = {30'd161, spc161_thread_id};

    wire[31:0] long_cpuid162;
    assign long_cpuid162 = {30'd162, spc162_thread_id};

    wire[31:0] long_cpuid163;
    assign long_cpuid163 = {30'd163, spc163_thread_id};

    wire[31:0] long_cpuid164;
    assign long_cpuid164 = {30'd164, spc164_thread_id};

    wire[31:0] long_cpuid165;
    assign long_cpuid165 = {30'd165, spc165_thread_id};

    wire[31:0] long_cpuid166;
    assign long_cpuid166 = {30'd166, spc166_thread_id};

    wire[31:0] long_cpuid167;
    assign long_cpuid167 = {30'd167, spc167_thread_id};

    wire[31:0] long_cpuid168;
    assign long_cpuid168 = {30'd168, spc168_thread_id};

    wire[31:0] long_cpuid169;
    assign long_cpuid169 = {30'd169, spc169_thread_id};

    wire[31:0] long_cpuid170;
    assign long_cpuid170 = {30'd170, spc170_thread_id};

    wire[31:0] long_cpuid171;
    assign long_cpuid171 = {30'd171, spc171_thread_id};

    wire[31:0] long_cpuid172;
    assign long_cpuid172 = {30'd172, spc172_thread_id};

    wire[31:0] long_cpuid173;
    assign long_cpuid173 = {30'd173, spc173_thread_id};

    wire[31:0] long_cpuid174;
    assign long_cpuid174 = {30'd174, spc174_thread_id};

    wire[31:0] long_cpuid175;
    assign long_cpuid175 = {30'd175, spc175_thread_id};

    wire[31:0] long_cpuid176;
    assign long_cpuid176 = {30'd176, spc176_thread_id};

    wire[31:0] long_cpuid177;
    assign long_cpuid177 = {30'd177, spc177_thread_id};

    wire[31:0] long_cpuid178;
    assign long_cpuid178 = {30'd178, spc178_thread_id};

    wire[31:0] long_cpuid179;
    assign long_cpuid179 = {30'd179, spc179_thread_id};

    wire[31:0] long_cpuid180;
    assign long_cpuid180 = {30'd180, spc180_thread_id};

    wire[31:0] long_cpuid181;
    assign long_cpuid181 = {30'd181, spc181_thread_id};

    wire[31:0] long_cpuid182;
    assign long_cpuid182 = {30'd182, spc182_thread_id};

    wire[31:0] long_cpuid183;
    assign long_cpuid183 = {30'd183, spc183_thread_id};

    wire[31:0] long_cpuid184;
    assign long_cpuid184 = {30'd184, spc184_thread_id};

    wire[31:0] long_cpuid185;
    assign long_cpuid185 = {30'd185, spc185_thread_id};

    wire[31:0] long_cpuid186;
    assign long_cpuid186 = {30'd186, spc186_thread_id};

    wire[31:0] long_cpuid187;
    assign long_cpuid187 = {30'd187, spc187_thread_id};

    wire[31:0] long_cpuid188;
    assign long_cpuid188 = {30'd188, spc188_thread_id};

    wire[31:0] long_cpuid189;
    assign long_cpuid189 = {30'd189, spc189_thread_id};

    wire[31:0] long_cpuid190;
    assign long_cpuid190 = {30'd190, spc190_thread_id};

    wire[31:0] long_cpuid191;
    assign long_cpuid191 = {30'd191, spc191_thread_id};

    wire[31:0] long_cpuid192;
    assign long_cpuid192 = {30'd192, spc192_thread_id};

    wire[31:0] long_cpuid193;
    assign long_cpuid193 = {30'd193, spc193_thread_id};

    wire[31:0] long_cpuid194;
    assign long_cpuid194 = {30'd194, spc194_thread_id};

    wire[31:0] long_cpuid195;
    assign long_cpuid195 = {30'd195, spc195_thread_id};

    wire[31:0] long_cpuid196;
    assign long_cpuid196 = {30'd196, spc196_thread_id};

    wire[31:0] long_cpuid197;
    assign long_cpuid197 = {30'd197, spc197_thread_id};

    wire[31:0] long_cpuid198;
    assign long_cpuid198 = {30'd198, spc198_thread_id};

    wire[31:0] long_cpuid199;
    assign long_cpuid199 = {30'd199, spc199_thread_id};

    wire[31:0] long_cpuid200;
    assign long_cpuid200 = {30'd200, spc200_thread_id};

    wire[31:0] long_cpuid201;
    assign long_cpuid201 = {30'd201, spc201_thread_id};

    wire[31:0] long_cpuid202;
    assign long_cpuid202 = {30'd202, spc202_thread_id};

    wire[31:0] long_cpuid203;
    assign long_cpuid203 = {30'd203, spc203_thread_id};

    wire[31:0] long_cpuid204;
    assign long_cpuid204 = {30'd204, spc204_thread_id};

    wire[31:0] long_cpuid205;
    assign long_cpuid205 = {30'd205, spc205_thread_id};

    wire[31:0] long_cpuid206;
    assign long_cpuid206 = {30'd206, spc206_thread_id};

    wire[31:0] long_cpuid207;
    assign long_cpuid207 = {30'd207, spc207_thread_id};

    wire[31:0] long_cpuid208;
    assign long_cpuid208 = {30'd208, spc208_thread_id};

    wire[31:0] long_cpuid209;
    assign long_cpuid209 = {30'd209, spc209_thread_id};

    wire[31:0] long_cpuid210;
    assign long_cpuid210 = {30'd210, spc210_thread_id};

    wire[31:0] long_cpuid211;
    assign long_cpuid211 = {30'd211, spc211_thread_id};

    wire[31:0] long_cpuid212;
    assign long_cpuid212 = {30'd212, spc212_thread_id};

    wire[31:0] long_cpuid213;
    assign long_cpuid213 = {30'd213, spc213_thread_id};

    wire[31:0] long_cpuid214;
    assign long_cpuid214 = {30'd214, spc214_thread_id};

    wire[31:0] long_cpuid215;
    assign long_cpuid215 = {30'd215, spc215_thread_id};

    wire[31:0] long_cpuid216;
    assign long_cpuid216 = {30'd216, spc216_thread_id};

    wire[31:0] long_cpuid217;
    assign long_cpuid217 = {30'd217, spc217_thread_id};

    wire[31:0] long_cpuid218;
    assign long_cpuid218 = {30'd218, spc218_thread_id};

    wire[31:0] long_cpuid219;
    assign long_cpuid219 = {30'd219, spc219_thread_id};

    wire[31:0] long_cpuid220;
    assign long_cpuid220 = {30'd220, spc220_thread_id};

    wire[31:0] long_cpuid221;
    assign long_cpuid221 = {30'd221, spc221_thread_id};

    wire[31:0] long_cpuid222;
    assign long_cpuid222 = {30'd222, spc222_thread_id};

    wire[31:0] long_cpuid223;
    assign long_cpuid223 = {30'd223, spc223_thread_id};

    wire[31:0] long_cpuid224;
    assign long_cpuid224 = {30'd224, spc224_thread_id};

    wire[31:0] long_cpuid225;
    assign long_cpuid225 = {30'd225, spc225_thread_id};

    wire[31:0] long_cpuid226;
    assign long_cpuid226 = {30'd226, spc226_thread_id};

    wire[31:0] long_cpuid227;
    assign long_cpuid227 = {30'd227, spc227_thread_id};

    wire[31:0] long_cpuid228;
    assign long_cpuid228 = {30'd228, spc228_thread_id};

    wire[31:0] long_cpuid229;
    assign long_cpuid229 = {30'd229, spc229_thread_id};

    wire[31:0] long_cpuid230;
    assign long_cpuid230 = {30'd230, spc230_thread_id};

    wire[31:0] long_cpuid231;
    assign long_cpuid231 = {30'd231, spc231_thread_id};

    wire[31:0] long_cpuid232;
    assign long_cpuid232 = {30'd232, spc232_thread_id};

    wire[31:0] long_cpuid233;
    assign long_cpuid233 = {30'd233, spc233_thread_id};

    wire[31:0] long_cpuid234;
    assign long_cpuid234 = {30'd234, spc234_thread_id};

    wire[31:0] long_cpuid235;
    assign long_cpuid235 = {30'd235, spc235_thread_id};

    wire[31:0] long_cpuid236;
    assign long_cpuid236 = {30'd236, spc236_thread_id};

    wire[31:0] long_cpuid237;
    assign long_cpuid237 = {30'd237, spc237_thread_id};

    wire[31:0] long_cpuid238;
    assign long_cpuid238 = {30'd238, spc238_thread_id};

    wire[31:0] long_cpuid239;
    assign long_cpuid239 = {30'd239, spc239_thread_id};

    wire[31:0] long_cpuid240;
    assign long_cpuid240 = {30'd240, spc240_thread_id};

    wire[31:0] long_cpuid241;
    assign long_cpuid241 = {30'd241, spc241_thread_id};

    wire[31:0] long_cpuid242;
    assign long_cpuid242 = {30'd242, spc242_thread_id};

    wire[31:0] long_cpuid243;
    assign long_cpuid243 = {30'd243, spc243_thread_id};

    wire[31:0] long_cpuid244;
    assign long_cpuid244 = {30'd244, spc244_thread_id};

    wire[31:0] long_cpuid245;
    assign long_cpuid245 = {30'd245, spc245_thread_id};

    wire[31:0] long_cpuid246;
    assign long_cpuid246 = {30'd246, spc246_thread_id};

    wire[31:0] long_cpuid247;
    assign long_cpuid247 = {30'd247, spc247_thread_id};

    wire[31:0] long_cpuid248;
    assign long_cpuid248 = {30'd248, spc248_thread_id};

    wire[31:0] long_cpuid249;
    assign long_cpuid249 = {30'd249, spc249_thread_id};

    wire[31:0] long_cpuid250;
    assign long_cpuid250 = {30'd250, spc250_thread_id};

    wire[31:0] long_cpuid251;
    assign long_cpuid251 = {30'd251, spc251_thread_id};

    wire[31:0] long_cpuid252;
    assign long_cpuid252 = {30'd252, spc252_thread_id};

    wire[31:0] long_cpuid253;
    assign long_cpuid253 = {30'd253, spc253_thread_id};

    wire[31:0] long_cpuid254;
    assign long_cpuid254 = {30'd254, spc254_thread_id};

    wire[31:0] long_cpuid255;
    assign long_cpuid255 = {30'd255, spc255_thread_id};

    wire[31:0] long_cpuid256;
    assign long_cpuid256 = {30'd256, spc256_thread_id};

    wire[31:0] long_cpuid257;
    assign long_cpuid257 = {30'd257, spc257_thread_id};

    wire[31:0] long_cpuid258;
    assign long_cpuid258 = {30'd258, spc258_thread_id};

    wire[31:0] long_cpuid259;
    assign long_cpuid259 = {30'd259, spc259_thread_id};

    wire[31:0] long_cpuid260;
    assign long_cpuid260 = {30'd260, spc260_thread_id};

    wire[31:0] long_cpuid261;
    assign long_cpuid261 = {30'd261, spc261_thread_id};

    wire[31:0] long_cpuid262;
    assign long_cpuid262 = {30'd262, spc262_thread_id};

    wire[31:0] long_cpuid263;
    assign long_cpuid263 = {30'd263, spc263_thread_id};

    wire[31:0] long_cpuid264;
    assign long_cpuid264 = {30'd264, spc264_thread_id};

    wire[31:0] long_cpuid265;
    assign long_cpuid265 = {30'd265, spc265_thread_id};

    wire[31:0] long_cpuid266;
    assign long_cpuid266 = {30'd266, spc266_thread_id};

    wire[31:0] long_cpuid267;
    assign long_cpuid267 = {30'd267, spc267_thread_id};

    wire[31:0] long_cpuid268;
    assign long_cpuid268 = {30'd268, spc268_thread_id};

    wire[31:0] long_cpuid269;
    assign long_cpuid269 = {30'd269, spc269_thread_id};

    wire[31:0] long_cpuid270;
    assign long_cpuid270 = {30'd270, spc270_thread_id};

    wire[31:0] long_cpuid271;
    assign long_cpuid271 = {30'd271, spc271_thread_id};

    wire[31:0] long_cpuid272;
    assign long_cpuid272 = {30'd272, spc272_thread_id};

    wire[31:0] long_cpuid273;
    assign long_cpuid273 = {30'd273, spc273_thread_id};

    wire[31:0] long_cpuid274;
    assign long_cpuid274 = {30'd274, spc274_thread_id};

    wire[31:0] long_cpuid275;
    assign long_cpuid275 = {30'd275, spc275_thread_id};

    wire[31:0] long_cpuid276;
    assign long_cpuid276 = {30'd276, spc276_thread_id};

    wire[31:0] long_cpuid277;
    assign long_cpuid277 = {30'd277, spc277_thread_id};

    wire[31:0] long_cpuid278;
    assign long_cpuid278 = {30'd278, spc278_thread_id};

    wire[31:0] long_cpuid279;
    assign long_cpuid279 = {30'd279, spc279_thread_id};

    wire[31:0] long_cpuid280;
    assign long_cpuid280 = {30'd280, spc280_thread_id};

    wire[31:0] long_cpuid281;
    assign long_cpuid281 = {30'd281, spc281_thread_id};

    wire[31:0] long_cpuid282;
    assign long_cpuid282 = {30'd282, spc282_thread_id};

    wire[31:0] long_cpuid283;
    assign long_cpuid283 = {30'd283, spc283_thread_id};

    wire[31:0] long_cpuid284;
    assign long_cpuid284 = {30'd284, spc284_thread_id};

    wire[31:0] long_cpuid285;
    assign long_cpuid285 = {30'd285, spc285_thread_id};

    wire[31:0] long_cpuid286;
    assign long_cpuid286 = {30'd286, spc286_thread_id};

    wire[31:0] long_cpuid287;
    assign long_cpuid287 = {30'd287, spc287_thread_id};

    wire[31:0] long_cpuid288;
    assign long_cpuid288 = {30'd288, spc288_thread_id};

    wire[31:0] long_cpuid289;
    assign long_cpuid289 = {30'd289, spc289_thread_id};

    wire[31:0] long_cpuid290;
    assign long_cpuid290 = {30'd290, spc290_thread_id};

    wire[31:0] long_cpuid291;
    assign long_cpuid291 = {30'd291, spc291_thread_id};

    wire[31:0] long_cpuid292;
    assign long_cpuid292 = {30'd292, spc292_thread_id};

    wire[31:0] long_cpuid293;
    assign long_cpuid293 = {30'd293, spc293_thread_id};

    wire[31:0] long_cpuid294;
    assign long_cpuid294 = {30'd294, spc294_thread_id};

    wire[31:0] long_cpuid295;
    assign long_cpuid295 = {30'd295, spc295_thread_id};

    wire[31:0] long_cpuid296;
    assign long_cpuid296 = {30'd296, spc296_thread_id};

    wire[31:0] long_cpuid297;
    assign long_cpuid297 = {30'd297, spc297_thread_id};

    wire[31:0] long_cpuid298;
    assign long_cpuid298 = {30'd298, spc298_thread_id};

    wire[31:0] long_cpuid299;
    assign long_cpuid299 = {30'd299, spc299_thread_id};

    wire[31:0] long_cpuid300;
    assign long_cpuid300 = {30'd300, spc300_thread_id};

    wire[31:0] long_cpuid301;
    assign long_cpuid301 = {30'd301, spc301_thread_id};

    wire[31:0] long_cpuid302;
    assign long_cpuid302 = {30'd302, spc302_thread_id};

    wire[31:0] long_cpuid303;
    assign long_cpuid303 = {30'd303, spc303_thread_id};

    wire[31:0] long_cpuid304;
    assign long_cpuid304 = {30'd304, spc304_thread_id};

    wire[31:0] long_cpuid305;
    assign long_cpuid305 = {30'd305, spc305_thread_id};

    wire[31:0] long_cpuid306;
    assign long_cpuid306 = {30'd306, spc306_thread_id};

    wire[31:0] long_cpuid307;
    assign long_cpuid307 = {30'd307, spc307_thread_id};

    wire[31:0] long_cpuid308;
    assign long_cpuid308 = {30'd308, spc308_thread_id};

    wire[31:0] long_cpuid309;
    assign long_cpuid309 = {30'd309, spc309_thread_id};

    wire[31:0] long_cpuid310;
    assign long_cpuid310 = {30'd310, spc310_thread_id};

    wire[31:0] long_cpuid311;
    assign long_cpuid311 = {30'd311, spc311_thread_id};

    wire[31:0] long_cpuid312;
    assign long_cpuid312 = {30'd312, spc312_thread_id};

    wire[31:0] long_cpuid313;
    assign long_cpuid313 = {30'd313, spc313_thread_id};

    wire[31:0] long_cpuid314;
    assign long_cpuid314 = {30'd314, spc314_thread_id};

    wire[31:0] long_cpuid315;
    assign long_cpuid315 = {30'd315, spc315_thread_id};

    wire[31:0] long_cpuid316;
    assign long_cpuid316 = {30'd316, spc316_thread_id};

    wire[31:0] long_cpuid317;
    assign long_cpuid317 = {30'd317, spc317_thread_id};

    wire[31:0] long_cpuid318;
    assign long_cpuid318 = {30'd318, spc318_thread_id};

    wire[31:0] long_cpuid319;
    assign long_cpuid319 = {30'd319, spc319_thread_id};

    wire[31:0] long_cpuid320;
    assign long_cpuid320 = {30'd320, spc320_thread_id};

    wire[31:0] long_cpuid321;
    assign long_cpuid321 = {30'd321, spc321_thread_id};

    wire[31:0] long_cpuid322;
    assign long_cpuid322 = {30'd322, spc322_thread_id};

    wire[31:0] long_cpuid323;
    assign long_cpuid323 = {30'd323, spc323_thread_id};

    wire[31:0] long_cpuid324;
    assign long_cpuid324 = {30'd324, spc324_thread_id};

    wire[31:0] long_cpuid325;
    assign long_cpuid325 = {30'd325, spc325_thread_id};

    wire[31:0] long_cpuid326;
    assign long_cpuid326 = {30'd326, spc326_thread_id};

    wire[31:0] long_cpuid327;
    assign long_cpuid327 = {30'd327, spc327_thread_id};

    wire[31:0] long_cpuid328;
    assign long_cpuid328 = {30'd328, spc328_thread_id};

    wire[31:0] long_cpuid329;
    assign long_cpuid329 = {30'd329, spc329_thread_id};

    wire[31:0] long_cpuid330;
    assign long_cpuid330 = {30'd330, spc330_thread_id};

    wire[31:0] long_cpuid331;
    assign long_cpuid331 = {30'd331, spc331_thread_id};

    wire[31:0] long_cpuid332;
    assign long_cpuid332 = {30'd332, spc332_thread_id};

    wire[31:0] long_cpuid333;
    assign long_cpuid333 = {30'd333, spc333_thread_id};

    wire[31:0] long_cpuid334;
    assign long_cpuid334 = {30'd334, spc334_thread_id};

    wire[31:0] long_cpuid335;
    assign long_cpuid335 = {30'd335, spc335_thread_id};

    wire[31:0] long_cpuid336;
    assign long_cpuid336 = {30'd336, spc336_thread_id};

    wire[31:0] long_cpuid337;
    assign long_cpuid337 = {30'd337, spc337_thread_id};

    wire[31:0] long_cpuid338;
    assign long_cpuid338 = {30'd338, spc338_thread_id};

    wire[31:0] long_cpuid339;
    assign long_cpuid339 = {30'd339, spc339_thread_id};

    wire[31:0] long_cpuid340;
    assign long_cpuid340 = {30'd340, spc340_thread_id};

    wire[31:0] long_cpuid341;
    assign long_cpuid341 = {30'd341, spc341_thread_id};

    wire[31:0] long_cpuid342;
    assign long_cpuid342 = {30'd342, spc342_thread_id};

    wire[31:0] long_cpuid343;
    assign long_cpuid343 = {30'd343, spc343_thread_id};

    wire[31:0] long_cpuid344;
    assign long_cpuid344 = {30'd344, spc344_thread_id};

    wire[31:0] long_cpuid345;
    assign long_cpuid345 = {30'd345, spc345_thread_id};

    wire[31:0] long_cpuid346;
    assign long_cpuid346 = {30'd346, spc346_thread_id};

    wire[31:0] long_cpuid347;
    assign long_cpuid347 = {30'd347, spc347_thread_id};

    wire[31:0] long_cpuid348;
    assign long_cpuid348 = {30'd348, spc348_thread_id};

    wire[31:0] long_cpuid349;
    assign long_cpuid349 = {30'd349, spc349_thread_id};

    wire[31:0] long_cpuid350;
    assign long_cpuid350 = {30'd350, spc350_thread_id};

    wire[31:0] long_cpuid351;
    assign long_cpuid351 = {30'd351, spc351_thread_id};

    wire[31:0] long_cpuid352;
    assign long_cpuid352 = {30'd352, spc352_thread_id};

    wire[31:0] long_cpuid353;
    assign long_cpuid353 = {30'd353, spc353_thread_id};

    wire[31:0] long_cpuid354;
    assign long_cpuid354 = {30'd354, spc354_thread_id};

    wire[31:0] long_cpuid355;
    assign long_cpuid355 = {30'd355, spc355_thread_id};

    wire[31:0] long_cpuid356;
    assign long_cpuid356 = {30'd356, spc356_thread_id};

    wire[31:0] long_cpuid357;
    assign long_cpuid357 = {30'd357, spc357_thread_id};

    wire[31:0] long_cpuid358;
    assign long_cpuid358 = {30'd358, spc358_thread_id};

    wire[31:0] long_cpuid359;
    assign long_cpuid359 = {30'd359, spc359_thread_id};

    wire[31:0] long_cpuid360;
    assign long_cpuid360 = {30'd360, spc360_thread_id};

    wire[31:0] long_cpuid361;
    assign long_cpuid361 = {30'd361, spc361_thread_id};

    wire[31:0] long_cpuid362;
    assign long_cpuid362 = {30'd362, spc362_thread_id};

    wire[31:0] long_cpuid363;
    assign long_cpuid363 = {30'd363, spc363_thread_id};

    wire[31:0] long_cpuid364;
    assign long_cpuid364 = {30'd364, spc364_thread_id};

    wire[31:0] long_cpuid365;
    assign long_cpuid365 = {30'd365, spc365_thread_id};

    wire[31:0] long_cpuid366;
    assign long_cpuid366 = {30'd366, spc366_thread_id};

    wire[31:0] long_cpuid367;
    assign long_cpuid367 = {30'd367, spc367_thread_id};

    wire[31:0] long_cpuid368;
    assign long_cpuid368 = {30'd368, spc368_thread_id};

    wire[31:0] long_cpuid369;
    assign long_cpuid369 = {30'd369, spc369_thread_id};

    wire[31:0] long_cpuid370;
    assign long_cpuid370 = {30'd370, spc370_thread_id};

    wire[31:0] long_cpuid371;
    assign long_cpuid371 = {30'd371, spc371_thread_id};

    wire[31:0] long_cpuid372;
    assign long_cpuid372 = {30'd372, spc372_thread_id};

    wire[31:0] long_cpuid373;
    assign long_cpuid373 = {30'd373, spc373_thread_id};

    wire[31:0] long_cpuid374;
    assign long_cpuid374 = {30'd374, spc374_thread_id};

    wire[31:0] long_cpuid375;
    assign long_cpuid375 = {30'd375, spc375_thread_id};

    wire[31:0] long_cpuid376;
    assign long_cpuid376 = {30'd376, spc376_thread_id};

    wire[31:0] long_cpuid377;
    assign long_cpuid377 = {30'd377, spc377_thread_id};

    wire[31:0] long_cpuid378;
    assign long_cpuid378 = {30'd378, spc378_thread_id};

    wire[31:0] long_cpuid379;
    assign long_cpuid379 = {30'd379, spc379_thread_id};

    wire[31:0] long_cpuid380;
    assign long_cpuid380 = {30'd380, spc380_thread_id};

    wire[31:0] long_cpuid381;
    assign long_cpuid381 = {30'd381, spc381_thread_id};

    wire[31:0] long_cpuid382;
    assign long_cpuid382 = {30'd382, spc382_thread_id};

    wire[31:0] long_cpuid383;
    assign long_cpuid383 = {30'd383, spc383_thread_id};

    wire[31:0] long_cpuid384;
    assign long_cpuid384 = {30'd384, spc384_thread_id};

    wire[31:0] long_cpuid385;
    assign long_cpuid385 = {30'd385, spc385_thread_id};

    wire[31:0] long_cpuid386;
    assign long_cpuid386 = {30'd386, spc386_thread_id};

    wire[31:0] long_cpuid387;
    assign long_cpuid387 = {30'd387, spc387_thread_id};

    wire[31:0] long_cpuid388;
    assign long_cpuid388 = {30'd388, spc388_thread_id};

    wire[31:0] long_cpuid389;
    assign long_cpuid389 = {30'd389, spc389_thread_id};

    wire[31:0] long_cpuid390;
    assign long_cpuid390 = {30'd390, spc390_thread_id};

    wire[31:0] long_cpuid391;
    assign long_cpuid391 = {30'd391, spc391_thread_id};

    wire[31:0] long_cpuid392;
    assign long_cpuid392 = {30'd392, spc392_thread_id};

    wire[31:0] long_cpuid393;
    assign long_cpuid393 = {30'd393, spc393_thread_id};

    wire[31:0] long_cpuid394;
    assign long_cpuid394 = {30'd394, spc394_thread_id};

    wire[31:0] long_cpuid395;
    assign long_cpuid395 = {30'd395, spc395_thread_id};

    wire[31:0] long_cpuid396;
    assign long_cpuid396 = {30'd396, spc396_thread_id};

    wire[31:0] long_cpuid397;
    assign long_cpuid397 = {30'd397, spc397_thread_id};

    wire[31:0] long_cpuid398;
    assign long_cpuid398 = {30'd398, spc398_thread_id};

    wire[31:0] long_cpuid399;
    assign long_cpuid399 = {30'd399, spc399_thread_id};

    wire[31:0] long_cpuid400;
    assign long_cpuid400 = {30'd400, spc400_thread_id};

    wire[31:0] long_cpuid401;
    assign long_cpuid401 = {30'd401, spc401_thread_id};

    wire[31:0] long_cpuid402;
    assign long_cpuid402 = {30'd402, spc402_thread_id};

    wire[31:0] long_cpuid403;
    assign long_cpuid403 = {30'd403, spc403_thread_id};

    wire[31:0] long_cpuid404;
    assign long_cpuid404 = {30'd404, spc404_thread_id};

    wire[31:0] long_cpuid405;
    assign long_cpuid405 = {30'd405, spc405_thread_id};

    wire[31:0] long_cpuid406;
    assign long_cpuid406 = {30'd406, spc406_thread_id};

    wire[31:0] long_cpuid407;
    assign long_cpuid407 = {30'd407, spc407_thread_id};

    wire[31:0] long_cpuid408;
    assign long_cpuid408 = {30'd408, spc408_thread_id};

    wire[31:0] long_cpuid409;
    assign long_cpuid409 = {30'd409, spc409_thread_id};

    wire[31:0] long_cpuid410;
    assign long_cpuid410 = {30'd410, spc410_thread_id};

    wire[31:0] long_cpuid411;
    assign long_cpuid411 = {30'd411, spc411_thread_id};

    wire[31:0] long_cpuid412;
    assign long_cpuid412 = {30'd412, spc412_thread_id};

    wire[31:0] long_cpuid413;
    assign long_cpuid413 = {30'd413, spc413_thread_id};

    wire[31:0] long_cpuid414;
    assign long_cpuid414 = {30'd414, spc414_thread_id};

    wire[31:0] long_cpuid415;
    assign long_cpuid415 = {30'd415, spc415_thread_id};

    wire[31:0] long_cpuid416;
    assign long_cpuid416 = {30'd416, spc416_thread_id};

    wire[31:0] long_cpuid417;
    assign long_cpuid417 = {30'd417, spc417_thread_id};

    wire[31:0] long_cpuid418;
    assign long_cpuid418 = {30'd418, spc418_thread_id};

    wire[31:0] long_cpuid419;
    assign long_cpuid419 = {30'd419, spc419_thread_id};

    wire[31:0] long_cpuid420;
    assign long_cpuid420 = {30'd420, spc420_thread_id};

    wire[31:0] long_cpuid421;
    assign long_cpuid421 = {30'd421, spc421_thread_id};

    wire[31:0] long_cpuid422;
    assign long_cpuid422 = {30'd422, spc422_thread_id};

    wire[31:0] long_cpuid423;
    assign long_cpuid423 = {30'd423, spc423_thread_id};

    wire[31:0] long_cpuid424;
    assign long_cpuid424 = {30'd424, spc424_thread_id};

    wire[31:0] long_cpuid425;
    assign long_cpuid425 = {30'd425, spc425_thread_id};

    wire[31:0] long_cpuid426;
    assign long_cpuid426 = {30'd426, spc426_thread_id};

    wire[31:0] long_cpuid427;
    assign long_cpuid427 = {30'd427, spc427_thread_id};

    wire[31:0] long_cpuid428;
    assign long_cpuid428 = {30'd428, spc428_thread_id};

    wire[31:0] long_cpuid429;
    assign long_cpuid429 = {30'd429, spc429_thread_id};

    wire[31:0] long_cpuid430;
    assign long_cpuid430 = {30'd430, spc430_thread_id};

    wire[31:0] long_cpuid431;
    assign long_cpuid431 = {30'd431, spc431_thread_id};

    wire[31:0] long_cpuid432;
    assign long_cpuid432 = {30'd432, spc432_thread_id};

    wire[31:0] long_cpuid433;
    assign long_cpuid433 = {30'd433, spc433_thread_id};

    wire[31:0] long_cpuid434;
    assign long_cpuid434 = {30'd434, spc434_thread_id};

    wire[31:0] long_cpuid435;
    assign long_cpuid435 = {30'd435, spc435_thread_id};

    wire[31:0] long_cpuid436;
    assign long_cpuid436 = {30'd436, spc436_thread_id};

    wire[31:0] long_cpuid437;
    assign long_cpuid437 = {30'd437, spc437_thread_id};

    wire[31:0] long_cpuid438;
    assign long_cpuid438 = {30'd438, spc438_thread_id};

    wire[31:0] long_cpuid439;
    assign long_cpuid439 = {30'd439, spc439_thread_id};

    wire[31:0] long_cpuid440;
    assign long_cpuid440 = {30'd440, spc440_thread_id};

    wire[31:0] long_cpuid441;
    assign long_cpuid441 = {30'd441, spc441_thread_id};

    wire[31:0] long_cpuid442;
    assign long_cpuid442 = {30'd442, spc442_thread_id};

    wire[31:0] long_cpuid443;
    assign long_cpuid443 = {30'd443, spc443_thread_id};

    wire[31:0] long_cpuid444;
    assign long_cpuid444 = {30'd444, spc444_thread_id};

    wire[31:0] long_cpuid445;
    assign long_cpuid445 = {30'd445, spc445_thread_id};

    wire[31:0] long_cpuid446;
    assign long_cpuid446 = {30'd446, spc446_thread_id};

    wire[31:0] long_cpuid447;
    assign long_cpuid447 = {30'd447, spc447_thread_id};

    wire[31:0] long_cpuid448;
    assign long_cpuid448 = {30'd448, spc448_thread_id};

    wire[31:0] long_cpuid449;
    assign long_cpuid449 = {30'd449, spc449_thread_id};

    wire[31:0] long_cpuid450;
    assign long_cpuid450 = {30'd450, spc450_thread_id};

    wire[31:0] long_cpuid451;
    assign long_cpuid451 = {30'd451, spc451_thread_id};

    wire[31:0] long_cpuid452;
    assign long_cpuid452 = {30'd452, spc452_thread_id};

    wire[31:0] long_cpuid453;
    assign long_cpuid453 = {30'd453, spc453_thread_id};

    wire[31:0] long_cpuid454;
    assign long_cpuid454 = {30'd454, spc454_thread_id};

    wire[31:0] long_cpuid455;
    assign long_cpuid455 = {30'd455, spc455_thread_id};

    wire[31:0] long_cpuid456;
    assign long_cpuid456 = {30'd456, spc456_thread_id};

    wire[31:0] long_cpuid457;
    assign long_cpuid457 = {30'd457, spc457_thread_id};

    wire[31:0] long_cpuid458;
    assign long_cpuid458 = {30'd458, spc458_thread_id};

    wire[31:0] long_cpuid459;
    assign long_cpuid459 = {30'd459, spc459_thread_id};

    wire[31:0] long_cpuid460;
    assign long_cpuid460 = {30'd460, spc460_thread_id};

    wire[31:0] long_cpuid461;
    assign long_cpuid461 = {30'd461, spc461_thread_id};

    wire[31:0] long_cpuid462;
    assign long_cpuid462 = {30'd462, spc462_thread_id};

    wire[31:0] long_cpuid463;
    assign long_cpuid463 = {30'd463, spc463_thread_id};

    wire[31:0] long_cpuid464;
    assign long_cpuid464 = {30'd464, spc464_thread_id};

    wire[31:0] long_cpuid465;
    assign long_cpuid465 = {30'd465, spc465_thread_id};

    wire[31:0] long_cpuid466;
    assign long_cpuid466 = {30'd466, spc466_thread_id};

    wire[31:0] long_cpuid467;
    assign long_cpuid467 = {30'd467, spc467_thread_id};

    wire[31:0] long_cpuid468;
    assign long_cpuid468 = {30'd468, spc468_thread_id};

    wire[31:0] long_cpuid469;
    assign long_cpuid469 = {30'd469, spc469_thread_id};

    wire[31:0] long_cpuid470;
    assign long_cpuid470 = {30'd470, spc470_thread_id};

    wire[31:0] long_cpuid471;
    assign long_cpuid471 = {30'd471, spc471_thread_id};

    wire[31:0] long_cpuid472;
    assign long_cpuid472 = {30'd472, spc472_thread_id};

    wire[31:0] long_cpuid473;
    assign long_cpuid473 = {30'd473, spc473_thread_id};

    wire[31:0] long_cpuid474;
    assign long_cpuid474 = {30'd474, spc474_thread_id};

    wire[31:0] long_cpuid475;
    assign long_cpuid475 = {30'd475, spc475_thread_id};

    wire[31:0] long_cpuid476;
    assign long_cpuid476 = {30'd476, spc476_thread_id};

    wire[31:0] long_cpuid477;
    assign long_cpuid477 = {30'd477, spc477_thread_id};

    wire[31:0] long_cpuid478;
    assign long_cpuid478 = {30'd478, spc478_thread_id};

    wire[31:0] long_cpuid479;
    assign long_cpuid479 = {30'd479, spc479_thread_id};

    wire[31:0] long_cpuid480;
    assign long_cpuid480 = {30'd480, spc480_thread_id};

    wire[31:0] long_cpuid481;
    assign long_cpuid481 = {30'd481, spc481_thread_id};

    wire[31:0] long_cpuid482;
    assign long_cpuid482 = {30'd482, spc482_thread_id};

    wire[31:0] long_cpuid483;
    assign long_cpuid483 = {30'd483, spc483_thread_id};

    wire[31:0] long_cpuid484;
    assign long_cpuid484 = {30'd484, spc484_thread_id};

    wire[31:0] long_cpuid485;
    assign long_cpuid485 = {30'd485, spc485_thread_id};

    wire[31:0] long_cpuid486;
    assign long_cpuid486 = {30'd486, spc486_thread_id};

    wire[31:0] long_cpuid487;
    assign long_cpuid487 = {30'd487, spc487_thread_id};

    wire[31:0] long_cpuid488;
    assign long_cpuid488 = {30'd488, spc488_thread_id};

    wire[31:0] long_cpuid489;
    assign long_cpuid489 = {30'd489, spc489_thread_id};

    wire[31:0] long_cpuid490;
    assign long_cpuid490 = {30'd490, spc490_thread_id};

    wire[31:0] long_cpuid491;
    assign long_cpuid491 = {30'd491, spc491_thread_id};

    wire[31:0] long_cpuid492;
    assign long_cpuid492 = {30'd492, spc492_thread_id};

    wire[31:0] long_cpuid493;
    assign long_cpuid493 = {30'd493, spc493_thread_id};

    wire[31:0] long_cpuid494;
    assign long_cpuid494 = {30'd494, spc494_thread_id};

    wire[31:0] long_cpuid495;
    assign long_cpuid495 = {30'd495, spc495_thread_id};

    wire[31:0] long_cpuid496;
    assign long_cpuid496 = {30'd496, spc496_thread_id};

    wire[31:0] long_cpuid497;
    assign long_cpuid497 = {30'd497, spc497_thread_id};

    wire[31:0] long_cpuid498;
    assign long_cpuid498 = {30'd498, spc498_thread_id};

    wire[31:0] long_cpuid499;
    assign long_cpuid499 = {30'd499, spc499_thread_id};

    wire[31:0] long_cpuid500;
    assign long_cpuid500 = {30'd500, spc500_thread_id};

    wire[31:0] long_cpuid501;
    assign long_cpuid501 = {30'd501, spc501_thread_id};

    wire[31:0] long_cpuid502;
    assign long_cpuid502 = {30'd502, spc502_thread_id};

    wire[31:0] long_cpuid503;
    assign long_cpuid503 = {30'd503, spc503_thread_id};

    wire[31:0] long_cpuid504;
    assign long_cpuid504 = {30'd504, spc504_thread_id};

    wire[31:0] long_cpuid505;
    assign long_cpuid505 = {30'd505, spc505_thread_id};

    wire[31:0] long_cpuid506;
    assign long_cpuid506 = {30'd506, spc506_thread_id};

    wire[31:0] long_cpuid507;
    assign long_cpuid507 = {30'd507, spc507_thread_id};

    wire[31:0] long_cpuid508;
    assign long_cpuid508 = {30'd508, spc508_thread_id};

    wire[31:0] long_cpuid509;
    assign long_cpuid509 = {30'd509, spc509_thread_id};

    wire[31:0] long_cpuid510;
    assign long_cpuid510 = {30'd510, spc510_thread_id};

    wire[31:0] long_cpuid511;
    assign long_cpuid511 = {30'd511, spc511_thread_id};

    wire[31:0] long_cpuid512;
    assign long_cpuid512 = {30'd512, spc512_thread_id};

    wire[31:0] long_cpuid513;
    assign long_cpuid513 = {30'd513, spc513_thread_id};

    wire[31:0] long_cpuid514;
    assign long_cpuid514 = {30'd514, spc514_thread_id};

    wire[31:0] long_cpuid515;
    assign long_cpuid515 = {30'd515, spc515_thread_id};

    wire[31:0] long_cpuid516;
    assign long_cpuid516 = {30'd516, spc516_thread_id};

    wire[31:0] long_cpuid517;
    assign long_cpuid517 = {30'd517, spc517_thread_id};

    wire[31:0] long_cpuid518;
    assign long_cpuid518 = {30'd518, spc518_thread_id};

    wire[31:0] long_cpuid519;
    assign long_cpuid519 = {30'd519, spc519_thread_id};

    wire[31:0] long_cpuid520;
    assign long_cpuid520 = {30'd520, spc520_thread_id};

    wire[31:0] long_cpuid521;
    assign long_cpuid521 = {30'd521, spc521_thread_id};

    wire[31:0] long_cpuid522;
    assign long_cpuid522 = {30'd522, spc522_thread_id};

    wire[31:0] long_cpuid523;
    assign long_cpuid523 = {30'd523, spc523_thread_id};

    wire[31:0] long_cpuid524;
    assign long_cpuid524 = {30'd524, spc524_thread_id};

    wire[31:0] long_cpuid525;
    assign long_cpuid525 = {30'd525, spc525_thread_id};

    wire[31:0] long_cpuid526;
    assign long_cpuid526 = {30'd526, spc526_thread_id};

    wire[31:0] long_cpuid527;
    assign long_cpuid527 = {30'd527, spc527_thread_id};

    wire[31:0] long_cpuid528;
    assign long_cpuid528 = {30'd528, spc528_thread_id};

    wire[31:0] long_cpuid529;
    assign long_cpuid529 = {30'd529, spc529_thread_id};

    wire[31:0] long_cpuid530;
    assign long_cpuid530 = {30'd530, spc530_thread_id};

    wire[31:0] long_cpuid531;
    assign long_cpuid531 = {30'd531, spc531_thread_id};

    wire[31:0] long_cpuid532;
    assign long_cpuid532 = {30'd532, spc532_thread_id};

    wire[31:0] long_cpuid533;
    assign long_cpuid533 = {30'd533, spc533_thread_id};

    wire[31:0] long_cpuid534;
    assign long_cpuid534 = {30'd534, spc534_thread_id};

    wire[31:0] long_cpuid535;
    assign long_cpuid535 = {30'd535, spc535_thread_id};

    wire[31:0] long_cpuid536;
    assign long_cpuid536 = {30'd536, spc536_thread_id};

    wire[31:0] long_cpuid537;
    assign long_cpuid537 = {30'd537, spc537_thread_id};

    wire[31:0] long_cpuid538;
    assign long_cpuid538 = {30'd538, spc538_thread_id};

    wire[31:0] long_cpuid539;
    assign long_cpuid539 = {30'd539, spc539_thread_id};

    wire[31:0] long_cpuid540;
    assign long_cpuid540 = {30'd540, spc540_thread_id};

    wire[31:0] long_cpuid541;
    assign long_cpuid541 = {30'd541, spc541_thread_id};

    wire[31:0] long_cpuid542;
    assign long_cpuid542 = {30'd542, spc542_thread_id};

    wire[31:0] long_cpuid543;
    assign long_cpuid543 = {30'd543, spc543_thread_id};

    wire[31:0] long_cpuid544;
    assign long_cpuid544 = {30'd544, spc544_thread_id};

    wire[31:0] long_cpuid545;
    assign long_cpuid545 = {30'd545, spc545_thread_id};

    wire[31:0] long_cpuid546;
    assign long_cpuid546 = {30'd546, spc546_thread_id};

    wire[31:0] long_cpuid547;
    assign long_cpuid547 = {30'd547, spc547_thread_id};

    wire[31:0] long_cpuid548;
    assign long_cpuid548 = {30'd548, spc548_thread_id};

    wire[31:0] long_cpuid549;
    assign long_cpuid549 = {30'd549, spc549_thread_id};

    wire[31:0] long_cpuid550;
    assign long_cpuid550 = {30'd550, spc550_thread_id};

    wire[31:0] long_cpuid551;
    assign long_cpuid551 = {30'd551, spc551_thread_id};

    wire[31:0] long_cpuid552;
    assign long_cpuid552 = {30'd552, spc552_thread_id};

    wire[31:0] long_cpuid553;
    assign long_cpuid553 = {30'd553, spc553_thread_id};

    wire[31:0] long_cpuid554;
    assign long_cpuid554 = {30'd554, spc554_thread_id};

    wire[31:0] long_cpuid555;
    assign long_cpuid555 = {30'd555, spc555_thread_id};

    wire[31:0] long_cpuid556;
    assign long_cpuid556 = {30'd556, spc556_thread_id};

    wire[31:0] long_cpuid557;
    assign long_cpuid557 = {30'd557, spc557_thread_id};

    wire[31:0] long_cpuid558;
    assign long_cpuid558 = {30'd558, spc558_thread_id};

    wire[31:0] long_cpuid559;
    assign long_cpuid559 = {30'd559, spc559_thread_id};

    wire[31:0] long_cpuid560;
    assign long_cpuid560 = {30'd560, spc560_thread_id};

    wire[31:0] long_cpuid561;
    assign long_cpuid561 = {30'd561, spc561_thread_id};

    wire[31:0] long_cpuid562;
    assign long_cpuid562 = {30'd562, spc562_thread_id};

    wire[31:0] long_cpuid563;
    assign long_cpuid563 = {30'd563, spc563_thread_id};

    wire[31:0] long_cpuid564;
    assign long_cpuid564 = {30'd564, spc564_thread_id};

    wire[31:0] long_cpuid565;
    assign long_cpuid565 = {30'd565, spc565_thread_id};

    wire[31:0] long_cpuid566;
    assign long_cpuid566 = {30'd566, spc566_thread_id};

    wire[31:0] long_cpuid567;
    assign long_cpuid567 = {30'd567, spc567_thread_id};

    wire[31:0] long_cpuid568;
    assign long_cpuid568 = {30'd568, spc568_thread_id};

    wire[31:0] long_cpuid569;
    assign long_cpuid569 = {30'd569, spc569_thread_id};

    wire[31:0] long_cpuid570;
    assign long_cpuid570 = {30'd570, spc570_thread_id};

    wire[31:0] long_cpuid571;
    assign long_cpuid571 = {30'd571, spc571_thread_id};

    wire[31:0] long_cpuid572;
    assign long_cpuid572 = {30'd572, spc572_thread_id};

    wire[31:0] long_cpuid573;
    assign long_cpuid573 = {30'd573, spc573_thread_id};

    wire[31:0] long_cpuid574;
    assign long_cpuid574 = {30'd574, spc574_thread_id};

    wire[31:0] long_cpuid575;
    assign long_cpuid575 = {30'd575, spc575_thread_id};

    wire[31:0] long_cpuid576;
    assign long_cpuid576 = {30'd576, spc576_thread_id};

    wire[31:0] long_cpuid577;
    assign long_cpuid577 = {30'd577, spc577_thread_id};

    wire[31:0] long_cpuid578;
    assign long_cpuid578 = {30'd578, spc578_thread_id};

    wire[31:0] long_cpuid579;
    assign long_cpuid579 = {30'd579, spc579_thread_id};

    wire[31:0] long_cpuid580;
    assign long_cpuid580 = {30'd580, spc580_thread_id};

    wire[31:0] long_cpuid581;
    assign long_cpuid581 = {30'd581, spc581_thread_id};

    wire[31:0] long_cpuid582;
    assign long_cpuid582 = {30'd582, spc582_thread_id};

    wire[31:0] long_cpuid583;
    assign long_cpuid583 = {30'd583, spc583_thread_id};

    wire[31:0] long_cpuid584;
    assign long_cpuid584 = {30'd584, spc584_thread_id};

    wire[31:0] long_cpuid585;
    assign long_cpuid585 = {30'd585, spc585_thread_id};

    wire[31:0] long_cpuid586;
    assign long_cpuid586 = {30'd586, spc586_thread_id};

    wire[31:0] long_cpuid587;
    assign long_cpuid587 = {30'd587, spc587_thread_id};

    wire[31:0] long_cpuid588;
    assign long_cpuid588 = {30'd588, spc588_thread_id};

    wire[31:0] long_cpuid589;
    assign long_cpuid589 = {30'd589, spc589_thread_id};

    wire[31:0] long_cpuid590;
    assign long_cpuid590 = {30'd590, spc590_thread_id};

    wire[31:0] long_cpuid591;
    assign long_cpuid591 = {30'd591, spc591_thread_id};

    wire[31:0] long_cpuid592;
    assign long_cpuid592 = {30'd592, spc592_thread_id};

    wire[31:0] long_cpuid593;
    assign long_cpuid593 = {30'd593, spc593_thread_id};

    wire[31:0] long_cpuid594;
    assign long_cpuid594 = {30'd594, spc594_thread_id};

    wire[31:0] long_cpuid595;
    assign long_cpuid595 = {30'd595, spc595_thread_id};

    wire[31:0] long_cpuid596;
    assign long_cpuid596 = {30'd596, spc596_thread_id};

    wire[31:0] long_cpuid597;
    assign long_cpuid597 = {30'd597, spc597_thread_id};

    wire[31:0] long_cpuid598;
    assign long_cpuid598 = {30'd598, spc598_thread_id};

    wire[31:0] long_cpuid599;
    assign long_cpuid599 = {30'd599, spc599_thread_id};

    wire[31:0] long_cpuid600;
    assign long_cpuid600 = {30'd600, spc600_thread_id};

    wire[31:0] long_cpuid601;
    assign long_cpuid601 = {30'd601, spc601_thread_id};

    wire[31:0] long_cpuid602;
    assign long_cpuid602 = {30'd602, spc602_thread_id};

    wire[31:0] long_cpuid603;
    assign long_cpuid603 = {30'd603, spc603_thread_id};

    wire[31:0] long_cpuid604;
    assign long_cpuid604 = {30'd604, spc604_thread_id};

    wire[31:0] long_cpuid605;
    assign long_cpuid605 = {30'd605, spc605_thread_id};

    wire[31:0] long_cpuid606;
    assign long_cpuid606 = {30'd606, spc606_thread_id};

    wire[31:0] long_cpuid607;
    assign long_cpuid607 = {30'd607, spc607_thread_id};

    wire[31:0] long_cpuid608;
    assign long_cpuid608 = {30'd608, spc608_thread_id};

    wire[31:0] long_cpuid609;
    assign long_cpuid609 = {30'd609, spc609_thread_id};

    wire[31:0] long_cpuid610;
    assign long_cpuid610 = {30'd610, spc610_thread_id};

    wire[31:0] long_cpuid611;
    assign long_cpuid611 = {30'd611, spc611_thread_id};

    wire[31:0] long_cpuid612;
    assign long_cpuid612 = {30'd612, spc612_thread_id};

    wire[31:0] long_cpuid613;
    assign long_cpuid613 = {30'd613, spc613_thread_id};

    wire[31:0] long_cpuid614;
    assign long_cpuid614 = {30'd614, spc614_thread_id};

    wire[31:0] long_cpuid615;
    assign long_cpuid615 = {30'd615, spc615_thread_id};

    wire[31:0] long_cpuid616;
    assign long_cpuid616 = {30'd616, spc616_thread_id};

    wire[31:0] long_cpuid617;
    assign long_cpuid617 = {30'd617, spc617_thread_id};

    wire[31:0] long_cpuid618;
    assign long_cpuid618 = {30'd618, spc618_thread_id};

    wire[31:0] long_cpuid619;
    assign long_cpuid619 = {30'd619, spc619_thread_id};

    wire[31:0] long_cpuid620;
    assign long_cpuid620 = {30'd620, spc620_thread_id};

    wire[31:0] long_cpuid621;
    assign long_cpuid621 = {30'd621, spc621_thread_id};

    wire[31:0] long_cpuid622;
    assign long_cpuid622 = {30'd622, spc622_thread_id};

    wire[31:0] long_cpuid623;
    assign long_cpuid623 = {30'd623, spc623_thread_id};

    wire[31:0] long_cpuid624;
    assign long_cpuid624 = {30'd624, spc624_thread_id};

    wire[31:0] long_cpuid625;
    assign long_cpuid625 = {30'd625, spc625_thread_id};

    wire[31:0] long_cpuid626;
    assign long_cpuid626 = {30'd626, spc626_thread_id};

    wire[31:0] long_cpuid627;
    assign long_cpuid627 = {30'd627, spc627_thread_id};

    wire[31:0] long_cpuid628;
    assign long_cpuid628 = {30'd628, spc628_thread_id};

    wire[31:0] long_cpuid629;
    assign long_cpuid629 = {30'd629, spc629_thread_id};

    wire[31:0] long_cpuid630;
    assign long_cpuid630 = {30'd630, spc630_thread_id};

    wire[31:0] long_cpuid631;
    assign long_cpuid631 = {30'd631, spc631_thread_id};

    wire[31:0] long_cpuid632;
    assign long_cpuid632 = {30'd632, spc632_thread_id};

    wire[31:0] long_cpuid633;
    assign long_cpuid633 = {30'd633, spc633_thread_id};

    wire[31:0] long_cpuid634;
    assign long_cpuid634 = {30'd634, spc634_thread_id};

    wire[31:0] long_cpuid635;
    assign long_cpuid635 = {30'd635, spc635_thread_id};

    wire[31:0] long_cpuid636;
    assign long_cpuid636 = {30'd636, spc636_thread_id};

    wire[31:0] long_cpuid637;
    assign long_cpuid637 = {30'd637, spc637_thread_id};

    wire[31:0] long_cpuid638;
    assign long_cpuid638 = {30'd638, spc638_thread_id};

    wire[31:0] long_cpuid639;
    assign long_cpuid639 = {30'd639, spc639_thread_id};

    wire[31:0] long_cpuid640;
    assign long_cpuid640 = {30'd640, spc640_thread_id};

    wire[31:0] long_cpuid641;
    assign long_cpuid641 = {30'd641, spc641_thread_id};

    wire[31:0] long_cpuid642;
    assign long_cpuid642 = {30'd642, spc642_thread_id};

    wire[31:0] long_cpuid643;
    assign long_cpuid643 = {30'd643, spc643_thread_id};

    wire[31:0] long_cpuid644;
    assign long_cpuid644 = {30'd644, spc644_thread_id};

    wire[31:0] long_cpuid645;
    assign long_cpuid645 = {30'd645, spc645_thread_id};

    wire[31:0] long_cpuid646;
    assign long_cpuid646 = {30'd646, spc646_thread_id};

    wire[31:0] long_cpuid647;
    assign long_cpuid647 = {30'd647, spc647_thread_id};

    wire[31:0] long_cpuid648;
    assign long_cpuid648 = {30'd648, spc648_thread_id};

    wire[31:0] long_cpuid649;
    assign long_cpuid649 = {30'd649, spc649_thread_id};

    wire[31:0] long_cpuid650;
    assign long_cpuid650 = {30'd650, spc650_thread_id};

    wire[31:0] long_cpuid651;
    assign long_cpuid651 = {30'd651, spc651_thread_id};

    wire[31:0] long_cpuid652;
    assign long_cpuid652 = {30'd652, spc652_thread_id};

    wire[31:0] long_cpuid653;
    assign long_cpuid653 = {30'd653, spc653_thread_id};

    wire[31:0] long_cpuid654;
    assign long_cpuid654 = {30'd654, spc654_thread_id};

    wire[31:0] long_cpuid655;
    assign long_cpuid655 = {30'd655, spc655_thread_id};

    wire[31:0] long_cpuid656;
    assign long_cpuid656 = {30'd656, spc656_thread_id};

    wire[31:0] long_cpuid657;
    assign long_cpuid657 = {30'd657, spc657_thread_id};

    wire[31:0] long_cpuid658;
    assign long_cpuid658 = {30'd658, spc658_thread_id};

    wire[31:0] long_cpuid659;
    assign long_cpuid659 = {30'd659, spc659_thread_id};

    wire[31:0] long_cpuid660;
    assign long_cpuid660 = {30'd660, spc660_thread_id};

    wire[31:0] long_cpuid661;
    assign long_cpuid661 = {30'd661, spc661_thread_id};

    wire[31:0] long_cpuid662;
    assign long_cpuid662 = {30'd662, spc662_thread_id};

    wire[31:0] long_cpuid663;
    assign long_cpuid663 = {30'd663, spc663_thread_id};

    wire[31:0] long_cpuid664;
    assign long_cpuid664 = {30'd664, spc664_thread_id};

    wire[31:0] long_cpuid665;
    assign long_cpuid665 = {30'd665, spc665_thread_id};

    wire[31:0] long_cpuid666;
    assign long_cpuid666 = {30'd666, spc666_thread_id};

    wire[31:0] long_cpuid667;
    assign long_cpuid667 = {30'd667, spc667_thread_id};

    wire[31:0] long_cpuid668;
    assign long_cpuid668 = {30'd668, spc668_thread_id};

    wire[31:0] long_cpuid669;
    assign long_cpuid669 = {30'd669, spc669_thread_id};

    wire[31:0] long_cpuid670;
    assign long_cpuid670 = {30'd670, spc670_thread_id};

    wire[31:0] long_cpuid671;
    assign long_cpuid671 = {30'd671, spc671_thread_id};

    wire[31:0] long_cpuid672;
    assign long_cpuid672 = {30'd672, spc672_thread_id};

    wire[31:0] long_cpuid673;
    assign long_cpuid673 = {30'd673, spc673_thread_id};

    wire[31:0] long_cpuid674;
    assign long_cpuid674 = {30'd674, spc674_thread_id};

    wire[31:0] long_cpuid675;
    assign long_cpuid675 = {30'd675, spc675_thread_id};

    wire[31:0] long_cpuid676;
    assign long_cpuid676 = {30'd676, spc676_thread_id};

    wire[31:0] long_cpuid677;
    assign long_cpuid677 = {30'd677, spc677_thread_id};

    wire[31:0] long_cpuid678;
    assign long_cpuid678 = {30'd678, spc678_thread_id};

    wire[31:0] long_cpuid679;
    assign long_cpuid679 = {30'd679, spc679_thread_id};

    wire[31:0] long_cpuid680;
    assign long_cpuid680 = {30'd680, spc680_thread_id};

    wire[31:0] long_cpuid681;
    assign long_cpuid681 = {30'd681, spc681_thread_id};

    wire[31:0] long_cpuid682;
    assign long_cpuid682 = {30'd682, spc682_thread_id};

    wire[31:0] long_cpuid683;
    assign long_cpuid683 = {30'd683, spc683_thread_id};

    wire[31:0] long_cpuid684;
    assign long_cpuid684 = {30'd684, spc684_thread_id};

    wire[31:0] long_cpuid685;
    assign long_cpuid685 = {30'd685, spc685_thread_id};

    wire[31:0] long_cpuid686;
    assign long_cpuid686 = {30'd686, spc686_thread_id};

    wire[31:0] long_cpuid687;
    assign long_cpuid687 = {30'd687, spc687_thread_id};

    wire[31:0] long_cpuid688;
    assign long_cpuid688 = {30'd688, spc688_thread_id};

    wire[31:0] long_cpuid689;
    assign long_cpuid689 = {30'd689, spc689_thread_id};

    wire[31:0] long_cpuid690;
    assign long_cpuid690 = {30'd690, spc690_thread_id};

    wire[31:0] long_cpuid691;
    assign long_cpuid691 = {30'd691, spc691_thread_id};

    wire[31:0] long_cpuid692;
    assign long_cpuid692 = {30'd692, spc692_thread_id};

    wire[31:0] long_cpuid693;
    assign long_cpuid693 = {30'd693, spc693_thread_id};

    wire[31:0] long_cpuid694;
    assign long_cpuid694 = {30'd694, spc694_thread_id};

    wire[31:0] long_cpuid695;
    assign long_cpuid695 = {30'd695, spc695_thread_id};

    wire[31:0] long_cpuid696;
    assign long_cpuid696 = {30'd696, spc696_thread_id};

    wire[31:0] long_cpuid697;
    assign long_cpuid697 = {30'd697, spc697_thread_id};

    wire[31:0] long_cpuid698;
    assign long_cpuid698 = {30'd698, spc698_thread_id};

    wire[31:0] long_cpuid699;
    assign long_cpuid699 = {30'd699, spc699_thread_id};

    wire[31:0] long_cpuid700;
    assign long_cpuid700 = {30'd700, spc700_thread_id};

    wire[31:0] long_cpuid701;
    assign long_cpuid701 = {30'd701, spc701_thread_id};

    wire[31:0] long_cpuid702;
    assign long_cpuid702 = {30'd702, spc702_thread_id};

    wire[31:0] long_cpuid703;
    assign long_cpuid703 = {30'd703, spc703_thread_id};

    wire[31:0] long_cpuid704;
    assign long_cpuid704 = {30'd704, spc704_thread_id};

    wire[31:0] long_cpuid705;
    assign long_cpuid705 = {30'd705, spc705_thread_id};

    wire[31:0] long_cpuid706;
    assign long_cpuid706 = {30'd706, spc706_thread_id};

    wire[31:0] long_cpuid707;
    assign long_cpuid707 = {30'd707, spc707_thread_id};

    wire[31:0] long_cpuid708;
    assign long_cpuid708 = {30'd708, spc708_thread_id};

    wire[31:0] long_cpuid709;
    assign long_cpuid709 = {30'd709, spc709_thread_id};

    wire[31:0] long_cpuid710;
    assign long_cpuid710 = {30'd710, spc710_thread_id};

    wire[31:0] long_cpuid711;
    assign long_cpuid711 = {30'd711, spc711_thread_id};

    wire[31:0] long_cpuid712;
    assign long_cpuid712 = {30'd712, spc712_thread_id};

    wire[31:0] long_cpuid713;
    assign long_cpuid713 = {30'd713, spc713_thread_id};

    wire[31:0] long_cpuid714;
    assign long_cpuid714 = {30'd714, spc714_thread_id};

    wire[31:0] long_cpuid715;
    assign long_cpuid715 = {30'd715, spc715_thread_id};

    wire[31:0] long_cpuid716;
    assign long_cpuid716 = {30'd716, spc716_thread_id};

    wire[31:0] long_cpuid717;
    assign long_cpuid717 = {30'd717, spc717_thread_id};

    wire[31:0] long_cpuid718;
    assign long_cpuid718 = {30'd718, spc718_thread_id};

    wire[31:0] long_cpuid719;
    assign long_cpuid719 = {30'd719, spc719_thread_id};

    wire[31:0] long_cpuid720;
    assign long_cpuid720 = {30'd720, spc720_thread_id};

    wire[31:0] long_cpuid721;
    assign long_cpuid721 = {30'd721, spc721_thread_id};

    wire[31:0] long_cpuid722;
    assign long_cpuid722 = {30'd722, spc722_thread_id};

    wire[31:0] long_cpuid723;
    assign long_cpuid723 = {30'd723, spc723_thread_id};

    wire[31:0] long_cpuid724;
    assign long_cpuid724 = {30'd724, spc724_thread_id};

    wire[31:0] long_cpuid725;
    assign long_cpuid725 = {30'd725, spc725_thread_id};

    wire[31:0] long_cpuid726;
    assign long_cpuid726 = {30'd726, spc726_thread_id};

    wire[31:0] long_cpuid727;
    assign long_cpuid727 = {30'd727, spc727_thread_id};

    wire[31:0] long_cpuid728;
    assign long_cpuid728 = {30'd728, spc728_thread_id};

    wire[31:0] long_cpuid729;
    assign long_cpuid729 = {30'd729, spc729_thread_id};

    wire[31:0] long_cpuid730;
    assign long_cpuid730 = {30'd730, spc730_thread_id};

    wire[31:0] long_cpuid731;
    assign long_cpuid731 = {30'd731, spc731_thread_id};

    wire[31:0] long_cpuid732;
    assign long_cpuid732 = {30'd732, spc732_thread_id};

    wire[31:0] long_cpuid733;
    assign long_cpuid733 = {30'd733, spc733_thread_id};

    wire[31:0] long_cpuid734;
    assign long_cpuid734 = {30'd734, spc734_thread_id};

    wire[31:0] long_cpuid735;
    assign long_cpuid735 = {30'd735, spc735_thread_id};

    wire[31:0] long_cpuid736;
    assign long_cpuid736 = {30'd736, spc736_thread_id};

    wire[31:0] long_cpuid737;
    assign long_cpuid737 = {30'd737, spc737_thread_id};

    wire[31:0] long_cpuid738;
    assign long_cpuid738 = {30'd738, spc738_thread_id};

    wire[31:0] long_cpuid739;
    assign long_cpuid739 = {30'd739, spc739_thread_id};

    wire[31:0] long_cpuid740;
    assign long_cpuid740 = {30'd740, spc740_thread_id};

    wire[31:0] long_cpuid741;
    assign long_cpuid741 = {30'd741, spc741_thread_id};

    wire[31:0] long_cpuid742;
    assign long_cpuid742 = {30'd742, spc742_thread_id};

    wire[31:0] long_cpuid743;
    assign long_cpuid743 = {30'd743, spc743_thread_id};

    wire[31:0] long_cpuid744;
    assign long_cpuid744 = {30'd744, spc744_thread_id};

    wire[31:0] long_cpuid745;
    assign long_cpuid745 = {30'd745, spc745_thread_id};

    wire[31:0] long_cpuid746;
    assign long_cpuid746 = {30'd746, spc746_thread_id};

    wire[31:0] long_cpuid747;
    assign long_cpuid747 = {30'd747, spc747_thread_id};

    wire[31:0] long_cpuid748;
    assign long_cpuid748 = {30'd748, spc748_thread_id};

    wire[31:0] long_cpuid749;
    assign long_cpuid749 = {30'd749, spc749_thread_id};

    wire[31:0] long_cpuid750;
    assign long_cpuid750 = {30'd750, spc750_thread_id};

    wire[31:0] long_cpuid751;
    assign long_cpuid751 = {30'd751, spc751_thread_id};

    wire[31:0] long_cpuid752;
    assign long_cpuid752 = {30'd752, spc752_thread_id};

    wire[31:0] long_cpuid753;
    assign long_cpuid753 = {30'd753, spc753_thread_id};

    wire[31:0] long_cpuid754;
    assign long_cpuid754 = {30'd754, spc754_thread_id};

    wire[31:0] long_cpuid755;
    assign long_cpuid755 = {30'd755, spc755_thread_id};

    wire[31:0] long_cpuid756;
    assign long_cpuid756 = {30'd756, spc756_thread_id};

    wire[31:0] long_cpuid757;
    assign long_cpuid757 = {30'd757, spc757_thread_id};

    wire[31:0] long_cpuid758;
    assign long_cpuid758 = {30'd758, spc758_thread_id};

    wire[31:0] long_cpuid759;
    assign long_cpuid759 = {30'd759, spc759_thread_id};

    wire[31:0] long_cpuid760;
    assign long_cpuid760 = {30'd760, spc760_thread_id};

    wire[31:0] long_cpuid761;
    assign long_cpuid761 = {30'd761, spc761_thread_id};

    wire[31:0] long_cpuid762;
    assign long_cpuid762 = {30'd762, spc762_thread_id};

    wire[31:0] long_cpuid763;
    assign long_cpuid763 = {30'd763, spc763_thread_id};

    wire[31:0] long_cpuid764;
    assign long_cpuid764 = {30'd764, spc764_thread_id};

    wire[31:0] long_cpuid765;
    assign long_cpuid765 = {30'd765, spc765_thread_id};

    wire[31:0] long_cpuid766;
    assign long_cpuid766 = {30'd766, spc766_thread_id};

    wire[31:0] long_cpuid767;
    assign long_cpuid767 = {30'd767, spc767_thread_id};

    wire[31:0] long_cpuid768;
    assign long_cpuid768 = {30'd768, spc768_thread_id};

    wire[31:0] long_cpuid769;
    assign long_cpuid769 = {30'd769, spc769_thread_id};

    wire[31:0] long_cpuid770;
    assign long_cpuid770 = {30'd770, spc770_thread_id};

    wire[31:0] long_cpuid771;
    assign long_cpuid771 = {30'd771, spc771_thread_id};

    wire[31:0] long_cpuid772;
    assign long_cpuid772 = {30'd772, spc772_thread_id};

    wire[31:0] long_cpuid773;
    assign long_cpuid773 = {30'd773, spc773_thread_id};

    wire[31:0] long_cpuid774;
    assign long_cpuid774 = {30'd774, spc774_thread_id};

    wire[31:0] long_cpuid775;
    assign long_cpuid775 = {30'd775, spc775_thread_id};

    wire[31:0] long_cpuid776;
    assign long_cpuid776 = {30'd776, spc776_thread_id};

    wire[31:0] long_cpuid777;
    assign long_cpuid777 = {30'd777, spc777_thread_id};

    wire[31:0] long_cpuid778;
    assign long_cpuid778 = {30'd778, spc778_thread_id};

    wire[31:0] long_cpuid779;
    assign long_cpuid779 = {30'd779, spc779_thread_id};

    wire[31:0] long_cpuid780;
    assign long_cpuid780 = {30'd780, spc780_thread_id};

    wire[31:0] long_cpuid781;
    assign long_cpuid781 = {30'd781, spc781_thread_id};

    wire[31:0] long_cpuid782;
    assign long_cpuid782 = {30'd782, spc782_thread_id};

    wire[31:0] long_cpuid783;
    assign long_cpuid783 = {30'd783, spc783_thread_id};

    wire[31:0] long_cpuid784;
    assign long_cpuid784 = {30'd784, spc784_thread_id};

    wire[31:0] long_cpuid785;
    assign long_cpuid785 = {30'd785, spc785_thread_id};

    wire[31:0] long_cpuid786;
    assign long_cpuid786 = {30'd786, spc786_thread_id};

    wire[31:0] long_cpuid787;
    assign long_cpuid787 = {30'd787, spc787_thread_id};

    wire[31:0] long_cpuid788;
    assign long_cpuid788 = {30'd788, spc788_thread_id};

    wire[31:0] long_cpuid789;
    assign long_cpuid789 = {30'd789, spc789_thread_id};

    wire[31:0] long_cpuid790;
    assign long_cpuid790 = {30'd790, spc790_thread_id};

    wire[31:0] long_cpuid791;
    assign long_cpuid791 = {30'd791, spc791_thread_id};

    wire[31:0] long_cpuid792;
    assign long_cpuid792 = {30'd792, spc792_thread_id};

    wire[31:0] long_cpuid793;
    assign long_cpuid793 = {30'd793, spc793_thread_id};

    wire[31:0] long_cpuid794;
    assign long_cpuid794 = {30'd794, spc794_thread_id};

    wire[31:0] long_cpuid795;
    assign long_cpuid795 = {30'd795, spc795_thread_id};

    wire[31:0] long_cpuid796;
    assign long_cpuid796 = {30'd796, spc796_thread_id};

    wire[31:0] long_cpuid797;
    assign long_cpuid797 = {30'd797, spc797_thread_id};

    wire[31:0] long_cpuid798;
    assign long_cpuid798 = {30'd798, spc798_thread_id};

    wire[31:0] long_cpuid799;
    assign long_cpuid799 = {30'd799, spc799_thread_id};

    wire[31:0] long_cpuid800;
    assign long_cpuid800 = {30'd800, spc800_thread_id};

    wire[31:0] long_cpuid801;
    assign long_cpuid801 = {30'd801, spc801_thread_id};

    wire[31:0] long_cpuid802;
    assign long_cpuid802 = {30'd802, spc802_thread_id};

    wire[31:0] long_cpuid803;
    assign long_cpuid803 = {30'd803, spc803_thread_id};

    wire[31:0] long_cpuid804;
    assign long_cpuid804 = {30'd804, spc804_thread_id};

    wire[31:0] long_cpuid805;
    assign long_cpuid805 = {30'd805, spc805_thread_id};

    wire[31:0] long_cpuid806;
    assign long_cpuid806 = {30'd806, spc806_thread_id};

    wire[31:0] long_cpuid807;
    assign long_cpuid807 = {30'd807, spc807_thread_id};

    wire[31:0] long_cpuid808;
    assign long_cpuid808 = {30'd808, spc808_thread_id};

    wire[31:0] long_cpuid809;
    assign long_cpuid809 = {30'd809, spc809_thread_id};

    wire[31:0] long_cpuid810;
    assign long_cpuid810 = {30'd810, spc810_thread_id};

    wire[31:0] long_cpuid811;
    assign long_cpuid811 = {30'd811, spc811_thread_id};

    wire[31:0] long_cpuid812;
    assign long_cpuid812 = {30'd812, spc812_thread_id};

    wire[31:0] long_cpuid813;
    assign long_cpuid813 = {30'd813, spc813_thread_id};

    wire[31:0] long_cpuid814;
    assign long_cpuid814 = {30'd814, spc814_thread_id};

    wire[31:0] long_cpuid815;
    assign long_cpuid815 = {30'd815, spc815_thread_id};

    wire[31:0] long_cpuid816;
    assign long_cpuid816 = {30'd816, spc816_thread_id};

    wire[31:0] long_cpuid817;
    assign long_cpuid817 = {30'd817, spc817_thread_id};

    wire[31:0] long_cpuid818;
    assign long_cpuid818 = {30'd818, spc818_thread_id};

    wire[31:0] long_cpuid819;
    assign long_cpuid819 = {30'd819, spc819_thread_id};

    wire[31:0] long_cpuid820;
    assign long_cpuid820 = {30'd820, spc820_thread_id};

    wire[31:0] long_cpuid821;
    assign long_cpuid821 = {30'd821, spc821_thread_id};

    wire[31:0] long_cpuid822;
    assign long_cpuid822 = {30'd822, spc822_thread_id};

    wire[31:0] long_cpuid823;
    assign long_cpuid823 = {30'd823, spc823_thread_id};

    wire[31:0] long_cpuid824;
    assign long_cpuid824 = {30'd824, spc824_thread_id};

    wire[31:0] long_cpuid825;
    assign long_cpuid825 = {30'd825, spc825_thread_id};

    wire[31:0] long_cpuid826;
    assign long_cpuid826 = {30'd826, spc826_thread_id};

    wire[31:0] long_cpuid827;
    assign long_cpuid827 = {30'd827, spc827_thread_id};

    wire[31:0] long_cpuid828;
    assign long_cpuid828 = {30'd828, spc828_thread_id};

    wire[31:0] long_cpuid829;
    assign long_cpuid829 = {30'd829, spc829_thread_id};

    wire[31:0] long_cpuid830;
    assign long_cpuid830 = {30'd830, spc830_thread_id};

    wire[31:0] long_cpuid831;
    assign long_cpuid831 = {30'd831, spc831_thread_id};

    wire[31:0] long_cpuid832;
    assign long_cpuid832 = {30'd832, spc832_thread_id};

    wire[31:0] long_cpuid833;
    assign long_cpuid833 = {30'd833, spc833_thread_id};

    wire[31:0] long_cpuid834;
    assign long_cpuid834 = {30'd834, spc834_thread_id};

    wire[31:0] long_cpuid835;
    assign long_cpuid835 = {30'd835, spc835_thread_id};

    wire[31:0] long_cpuid836;
    assign long_cpuid836 = {30'd836, spc836_thread_id};

    wire[31:0] long_cpuid837;
    assign long_cpuid837 = {30'd837, spc837_thread_id};

    wire[31:0] long_cpuid838;
    assign long_cpuid838 = {30'd838, spc838_thread_id};

    wire[31:0] long_cpuid839;
    assign long_cpuid839 = {30'd839, spc839_thread_id};

    wire[31:0] long_cpuid840;
    assign long_cpuid840 = {30'd840, spc840_thread_id};

    wire[31:0] long_cpuid841;
    assign long_cpuid841 = {30'd841, spc841_thread_id};

    wire[31:0] long_cpuid842;
    assign long_cpuid842 = {30'd842, spc842_thread_id};

    wire[31:0] long_cpuid843;
    assign long_cpuid843 = {30'd843, spc843_thread_id};

    wire[31:0] long_cpuid844;
    assign long_cpuid844 = {30'd844, spc844_thread_id};

    wire[31:0] long_cpuid845;
    assign long_cpuid845 = {30'd845, spc845_thread_id};

    wire[31:0] long_cpuid846;
    assign long_cpuid846 = {30'd846, spc846_thread_id};

    wire[31:0] long_cpuid847;
    assign long_cpuid847 = {30'd847, spc847_thread_id};

    wire[31:0] long_cpuid848;
    assign long_cpuid848 = {30'd848, spc848_thread_id};

    wire[31:0] long_cpuid849;
    assign long_cpuid849 = {30'd849, spc849_thread_id};

    wire[31:0] long_cpuid850;
    assign long_cpuid850 = {30'd850, spc850_thread_id};

    wire[31:0] long_cpuid851;
    assign long_cpuid851 = {30'd851, spc851_thread_id};

    wire[31:0] long_cpuid852;
    assign long_cpuid852 = {30'd852, spc852_thread_id};

    wire[31:0] long_cpuid853;
    assign long_cpuid853 = {30'd853, spc853_thread_id};

    wire[31:0] long_cpuid854;
    assign long_cpuid854 = {30'd854, spc854_thread_id};

    wire[31:0] long_cpuid855;
    assign long_cpuid855 = {30'd855, spc855_thread_id};

    wire[31:0] long_cpuid856;
    assign long_cpuid856 = {30'd856, spc856_thread_id};

    wire[31:0] long_cpuid857;
    assign long_cpuid857 = {30'd857, spc857_thread_id};

    wire[31:0] long_cpuid858;
    assign long_cpuid858 = {30'd858, spc858_thread_id};

    wire[31:0] long_cpuid859;
    assign long_cpuid859 = {30'd859, spc859_thread_id};

    wire[31:0] long_cpuid860;
    assign long_cpuid860 = {30'd860, spc860_thread_id};

    wire[31:0] long_cpuid861;
    assign long_cpuid861 = {30'd861, spc861_thread_id};

    wire[31:0] long_cpuid862;
    assign long_cpuid862 = {30'd862, spc862_thread_id};

    wire[31:0] long_cpuid863;
    assign long_cpuid863 = {30'd863, spc863_thread_id};

    wire[31:0] long_cpuid864;
    assign long_cpuid864 = {30'd864, spc864_thread_id};

    wire[31:0] long_cpuid865;
    assign long_cpuid865 = {30'd865, spc865_thread_id};

    wire[31:0] long_cpuid866;
    assign long_cpuid866 = {30'd866, spc866_thread_id};

    wire[31:0] long_cpuid867;
    assign long_cpuid867 = {30'd867, spc867_thread_id};

    wire[31:0] long_cpuid868;
    assign long_cpuid868 = {30'd868, spc868_thread_id};

    wire[31:0] long_cpuid869;
    assign long_cpuid869 = {30'd869, spc869_thread_id};

    wire[31:0] long_cpuid870;
    assign long_cpuid870 = {30'd870, spc870_thread_id};

    wire[31:0] long_cpuid871;
    assign long_cpuid871 = {30'd871, spc871_thread_id};

    wire[31:0] long_cpuid872;
    assign long_cpuid872 = {30'd872, spc872_thread_id};

    wire[31:0] long_cpuid873;
    assign long_cpuid873 = {30'd873, spc873_thread_id};

    wire[31:0] long_cpuid874;
    assign long_cpuid874 = {30'd874, spc874_thread_id};

    wire[31:0] long_cpuid875;
    assign long_cpuid875 = {30'd875, spc875_thread_id};

    wire[31:0] long_cpuid876;
    assign long_cpuid876 = {30'd876, spc876_thread_id};

    wire[31:0] long_cpuid877;
    assign long_cpuid877 = {30'd877, spc877_thread_id};

    wire[31:0] long_cpuid878;
    assign long_cpuid878 = {30'd878, spc878_thread_id};

    wire[31:0] long_cpuid879;
    assign long_cpuid879 = {30'd879, spc879_thread_id};

    wire[31:0] long_cpuid880;
    assign long_cpuid880 = {30'd880, spc880_thread_id};

    wire[31:0] long_cpuid881;
    assign long_cpuid881 = {30'd881, spc881_thread_id};

    wire[31:0] long_cpuid882;
    assign long_cpuid882 = {30'd882, spc882_thread_id};

    wire[31:0] long_cpuid883;
    assign long_cpuid883 = {30'd883, spc883_thread_id};

    wire[31:0] long_cpuid884;
    assign long_cpuid884 = {30'd884, spc884_thread_id};

    wire[31:0] long_cpuid885;
    assign long_cpuid885 = {30'd885, spc885_thread_id};

    wire[31:0] long_cpuid886;
    assign long_cpuid886 = {30'd886, spc886_thread_id};

    wire[31:0] long_cpuid887;
    assign long_cpuid887 = {30'd887, spc887_thread_id};

    wire[31:0] long_cpuid888;
    assign long_cpuid888 = {30'd888, spc888_thread_id};

    wire[31:0] long_cpuid889;
    assign long_cpuid889 = {30'd889, spc889_thread_id};

    wire[31:0] long_cpuid890;
    assign long_cpuid890 = {30'd890, spc890_thread_id};

    wire[31:0] long_cpuid891;
    assign long_cpuid891 = {30'd891, spc891_thread_id};

    wire[31:0] long_cpuid892;
    assign long_cpuid892 = {30'd892, spc892_thread_id};

    wire[31:0] long_cpuid893;
    assign long_cpuid893 = {30'd893, spc893_thread_id};

    wire[31:0] long_cpuid894;
    assign long_cpuid894 = {30'd894, spc894_thread_id};

    wire[31:0] long_cpuid895;
    assign long_cpuid895 = {30'd895, spc895_thread_id};

    wire[31:0] long_cpuid896;
    assign long_cpuid896 = {30'd896, spc896_thread_id};

    wire[31:0] long_cpuid897;
    assign long_cpuid897 = {30'd897, spc897_thread_id};

    wire[31:0] long_cpuid898;
    assign long_cpuid898 = {30'd898, spc898_thread_id};

    wire[31:0] long_cpuid899;
    assign long_cpuid899 = {30'd899, spc899_thread_id};

    wire[31:0] long_cpuid900;
    assign long_cpuid900 = {30'd900, spc900_thread_id};

    wire[31:0] long_cpuid901;
    assign long_cpuid901 = {30'd901, spc901_thread_id};

    wire[31:0] long_cpuid902;
    assign long_cpuid902 = {30'd902, spc902_thread_id};

    wire[31:0] long_cpuid903;
    assign long_cpuid903 = {30'd903, spc903_thread_id};

    wire[31:0] long_cpuid904;
    assign long_cpuid904 = {30'd904, spc904_thread_id};

    wire[31:0] long_cpuid905;
    assign long_cpuid905 = {30'd905, spc905_thread_id};

    wire[31:0] long_cpuid906;
    assign long_cpuid906 = {30'd906, spc906_thread_id};

    wire[31:0] long_cpuid907;
    assign long_cpuid907 = {30'd907, spc907_thread_id};

    wire[31:0] long_cpuid908;
    assign long_cpuid908 = {30'd908, spc908_thread_id};

    wire[31:0] long_cpuid909;
    assign long_cpuid909 = {30'd909, spc909_thread_id};

    wire[31:0] long_cpuid910;
    assign long_cpuid910 = {30'd910, spc910_thread_id};

    wire[31:0] long_cpuid911;
    assign long_cpuid911 = {30'd911, spc911_thread_id};

    wire[31:0] long_cpuid912;
    assign long_cpuid912 = {30'd912, spc912_thread_id};

    wire[31:0] long_cpuid913;
    assign long_cpuid913 = {30'd913, spc913_thread_id};

    wire[31:0] long_cpuid914;
    assign long_cpuid914 = {30'd914, spc914_thread_id};

    wire[31:0] long_cpuid915;
    assign long_cpuid915 = {30'd915, spc915_thread_id};

    wire[31:0] long_cpuid916;
    assign long_cpuid916 = {30'd916, spc916_thread_id};

    wire[31:0] long_cpuid917;
    assign long_cpuid917 = {30'd917, spc917_thread_id};

    wire[31:0] long_cpuid918;
    assign long_cpuid918 = {30'd918, spc918_thread_id};

    wire[31:0] long_cpuid919;
    assign long_cpuid919 = {30'd919, spc919_thread_id};

    wire[31:0] long_cpuid920;
    assign long_cpuid920 = {30'd920, spc920_thread_id};

    wire[31:0] long_cpuid921;
    assign long_cpuid921 = {30'd921, spc921_thread_id};

    wire[31:0] long_cpuid922;
    assign long_cpuid922 = {30'd922, spc922_thread_id};

    wire[31:0] long_cpuid923;
    assign long_cpuid923 = {30'd923, spc923_thread_id};

    wire[31:0] long_cpuid924;
    assign long_cpuid924 = {30'd924, spc924_thread_id};

    wire[31:0] long_cpuid925;
    assign long_cpuid925 = {30'd925, spc925_thread_id};

    wire[31:0] long_cpuid926;
    assign long_cpuid926 = {30'd926, spc926_thread_id};

    wire[31:0] long_cpuid927;
    assign long_cpuid927 = {30'd927, spc927_thread_id};

    wire[31:0] long_cpuid928;
    assign long_cpuid928 = {30'd928, spc928_thread_id};

    wire[31:0] long_cpuid929;
    assign long_cpuid929 = {30'd929, spc929_thread_id};

    wire[31:0] long_cpuid930;
    assign long_cpuid930 = {30'd930, spc930_thread_id};

    wire[31:0] long_cpuid931;
    assign long_cpuid931 = {30'd931, spc931_thread_id};

    wire[31:0] long_cpuid932;
    assign long_cpuid932 = {30'd932, spc932_thread_id};

    wire[31:0] long_cpuid933;
    assign long_cpuid933 = {30'd933, spc933_thread_id};

    wire[31:0] long_cpuid934;
    assign long_cpuid934 = {30'd934, spc934_thread_id};

    wire[31:0] long_cpuid935;
    assign long_cpuid935 = {30'd935, spc935_thread_id};

    wire[31:0] long_cpuid936;
    assign long_cpuid936 = {30'd936, spc936_thread_id};

    wire[31:0] long_cpuid937;
    assign long_cpuid937 = {30'd937, spc937_thread_id};

    wire[31:0] long_cpuid938;
    assign long_cpuid938 = {30'd938, spc938_thread_id};

    wire[31:0] long_cpuid939;
    assign long_cpuid939 = {30'd939, spc939_thread_id};

    wire[31:0] long_cpuid940;
    assign long_cpuid940 = {30'd940, spc940_thread_id};

    wire[31:0] long_cpuid941;
    assign long_cpuid941 = {30'd941, spc941_thread_id};

    wire[31:0] long_cpuid942;
    assign long_cpuid942 = {30'd942, spc942_thread_id};

    wire[31:0] long_cpuid943;
    assign long_cpuid943 = {30'd943, spc943_thread_id};

    wire[31:0] long_cpuid944;
    assign long_cpuid944 = {30'd944, spc944_thread_id};

    wire[31:0] long_cpuid945;
    assign long_cpuid945 = {30'd945, spc945_thread_id};

    wire[31:0] long_cpuid946;
    assign long_cpuid946 = {30'd946, spc946_thread_id};

    wire[31:0] long_cpuid947;
    assign long_cpuid947 = {30'd947, spc947_thread_id};

    wire[31:0] long_cpuid948;
    assign long_cpuid948 = {30'd948, spc948_thread_id};

    wire[31:0] long_cpuid949;
    assign long_cpuid949 = {30'd949, spc949_thread_id};

    wire[31:0] long_cpuid950;
    assign long_cpuid950 = {30'd950, spc950_thread_id};

    wire[31:0] long_cpuid951;
    assign long_cpuid951 = {30'd951, spc951_thread_id};

    wire[31:0] long_cpuid952;
    assign long_cpuid952 = {30'd952, spc952_thread_id};

    wire[31:0] long_cpuid953;
    assign long_cpuid953 = {30'd953, spc953_thread_id};

    wire[31:0] long_cpuid954;
    assign long_cpuid954 = {30'd954, spc954_thread_id};

    wire[31:0] long_cpuid955;
    assign long_cpuid955 = {30'd955, spc955_thread_id};

    wire[31:0] long_cpuid956;
    assign long_cpuid956 = {30'd956, spc956_thread_id};

    wire[31:0] long_cpuid957;
    assign long_cpuid957 = {30'd957, spc957_thread_id};

    wire[31:0] long_cpuid958;
    assign long_cpuid958 = {30'd958, spc958_thread_id};

    wire[31:0] long_cpuid959;
    assign long_cpuid959 = {30'd959, spc959_thread_id};

    wire[31:0] long_cpuid960;
    assign long_cpuid960 = {30'd960, spc960_thread_id};

    wire[31:0] long_cpuid961;
    assign long_cpuid961 = {30'd961, spc961_thread_id};

    wire[31:0] long_cpuid962;
    assign long_cpuid962 = {30'd962, spc962_thread_id};

    wire[31:0] long_cpuid963;
    assign long_cpuid963 = {30'd963, spc963_thread_id};

    wire[31:0] long_cpuid964;
    assign long_cpuid964 = {30'd964, spc964_thread_id};

    wire[31:0] long_cpuid965;
    assign long_cpuid965 = {30'd965, spc965_thread_id};

    wire[31:0] long_cpuid966;
    assign long_cpuid966 = {30'd966, spc966_thread_id};

    wire[31:0] long_cpuid967;
    assign long_cpuid967 = {30'd967, spc967_thread_id};

    wire[31:0] long_cpuid968;
    assign long_cpuid968 = {30'd968, spc968_thread_id};

    wire[31:0] long_cpuid969;
    assign long_cpuid969 = {30'd969, spc969_thread_id};

    wire[31:0] long_cpuid970;
    assign long_cpuid970 = {30'd970, spc970_thread_id};

    wire[31:0] long_cpuid971;
    assign long_cpuid971 = {30'd971, spc971_thread_id};

    wire[31:0] long_cpuid972;
    assign long_cpuid972 = {30'd972, spc972_thread_id};

    wire[31:0] long_cpuid973;
    assign long_cpuid973 = {30'd973, spc973_thread_id};

    wire[31:0] long_cpuid974;
    assign long_cpuid974 = {30'd974, spc974_thread_id};

    wire[31:0] long_cpuid975;
    assign long_cpuid975 = {30'd975, spc975_thread_id};

    wire[31:0] long_cpuid976;
    assign long_cpuid976 = {30'd976, spc976_thread_id};

    wire[31:0] long_cpuid977;
    assign long_cpuid977 = {30'd977, spc977_thread_id};

    wire[31:0] long_cpuid978;
    assign long_cpuid978 = {30'd978, spc978_thread_id};

    wire[31:0] long_cpuid979;
    assign long_cpuid979 = {30'd979, spc979_thread_id};

    wire[31:0] long_cpuid980;
    assign long_cpuid980 = {30'd980, spc980_thread_id};

    wire[31:0] long_cpuid981;
    assign long_cpuid981 = {30'd981, spc981_thread_id};

    wire[31:0] long_cpuid982;
    assign long_cpuid982 = {30'd982, spc982_thread_id};

    wire[31:0] long_cpuid983;
    assign long_cpuid983 = {30'd983, spc983_thread_id};

    wire[31:0] long_cpuid984;
    assign long_cpuid984 = {30'd984, spc984_thread_id};

    wire[31:0] long_cpuid985;
    assign long_cpuid985 = {30'd985, spc985_thread_id};

    wire[31:0] long_cpuid986;
    assign long_cpuid986 = {30'd986, spc986_thread_id};

    wire[31:0] long_cpuid987;
    assign long_cpuid987 = {30'd987, spc987_thread_id};

    wire[31:0] long_cpuid988;
    assign long_cpuid988 = {30'd988, spc988_thread_id};

    wire[31:0] long_cpuid989;
    assign long_cpuid989 = {30'd989, spc989_thread_id};

    wire[31:0] long_cpuid990;
    assign long_cpuid990 = {30'd990, spc990_thread_id};

    wire[31:0] long_cpuid991;
    assign long_cpuid991 = {30'd991, spc991_thread_id};

    wire[31:0] long_cpuid992;
    assign long_cpuid992 = {30'd992, spc992_thread_id};

    wire[31:0] long_cpuid993;
    assign long_cpuid993 = {30'd993, spc993_thread_id};

    wire[31:0] long_cpuid994;
    assign long_cpuid994 = {30'd994, spc994_thread_id};

    wire[31:0] long_cpuid995;
    assign long_cpuid995 = {30'd995, spc995_thread_id};

    wire[31:0] long_cpuid996;
    assign long_cpuid996 = {30'd996, spc996_thread_id};

    wire[31:0] long_cpuid997;
    assign long_cpuid997 = {30'd997, spc997_thread_id};

    wire[31:0] long_cpuid998;
    assign long_cpuid998 = {30'd998, spc998_thread_id};

    wire[31:0] long_cpuid999;
    assign long_cpuid999 = {30'd999, spc999_thread_id};

    wire[31:0] long_cpuid1000;
    assign long_cpuid1000 = {30'd1000, spc1000_thread_id};

    wire[31:0] long_cpuid1001;
    assign long_cpuid1001 = {30'd1001, spc1001_thread_id};

    wire[31:0] long_cpuid1002;
    assign long_cpuid1002 = {30'd1002, spc1002_thread_id};

    wire[31:0] long_cpuid1003;
    assign long_cpuid1003 = {30'd1003, spc1003_thread_id};

    wire[31:0] long_cpuid1004;
    assign long_cpuid1004 = {30'd1004, spc1004_thread_id};

    wire[31:0] long_cpuid1005;
    assign long_cpuid1005 = {30'd1005, spc1005_thread_id};

    wire[31:0] long_cpuid1006;
    assign long_cpuid1006 = {30'd1006, spc1006_thread_id};

    wire[31:0] long_cpuid1007;
    assign long_cpuid1007 = {30'd1007, spc1007_thread_id};

    wire[31:0] long_cpuid1008;
    assign long_cpuid1008 = {30'd1008, spc1008_thread_id};

    wire[31:0] long_cpuid1009;
    assign long_cpuid1009 = {30'd1009, spc1009_thread_id};

    wire[31:0] long_cpuid1010;
    assign long_cpuid1010 = {30'd1010, spc1010_thread_id};

    wire[31:0] long_cpuid1011;
    assign long_cpuid1011 = {30'd1011, spc1011_thread_id};

    wire[31:0] long_cpuid1012;
    assign long_cpuid1012 = {30'd1012, spc1012_thread_id};

    wire[31:0] long_cpuid1013;
    assign long_cpuid1013 = {30'd1013, spc1013_thread_id};

    wire[31:0] long_cpuid1014;
    assign long_cpuid1014 = {30'd1014, spc1014_thread_id};

    wire[31:0] long_cpuid1015;
    assign long_cpuid1015 = {30'd1015, spc1015_thread_id};

    wire[31:0] long_cpuid1016;
    assign long_cpuid1016 = {30'd1016, spc1016_thread_id};

    wire[31:0] long_cpuid1017;
    assign long_cpuid1017 = {30'd1017, spc1017_thread_id};

    wire[31:0] long_cpuid1018;
    assign long_cpuid1018 = {30'd1018, spc1018_thread_id};

    wire[31:0] long_cpuid1019;
    assign long_cpuid1019 = {30'd1019, spc1019_thread_id};

    wire[31:0] long_cpuid1020;
    assign long_cpuid1020 = {30'd1020, spc1020_thread_id};

    wire[31:0] long_cpuid1021;
    assign long_cpuid1021 = {30'd1021, spc1021_thread_id};

    wire[31:0] long_cpuid1022;
    assign long_cpuid1022 = {30'd1022, spc1022_thread_id};

    wire[31:0] long_cpuid1023;
    assign long_cpuid1023 = {30'd1023, spc1023_thread_id};


always @* begin
done[0]   = spc0_inst_done;//sparc 0
done[1]   = spc1_inst_done;//sparc 1
done[2]   = spc2_inst_done;//sparc 2
done[3]   = spc3_inst_done;//sparc 3
done[4]   = spc4_inst_done;//sparc 4
done[5]   = spc5_inst_done;//sparc 5
done[6]   = spc6_inst_done;//sparc 6
done[7]   = spc7_inst_done;//sparc 7
done[8]   = spc8_inst_done;//sparc 8
done[9]   = spc9_inst_done;//sparc 9
done[10]   = spc10_inst_done;//sparc 10
done[11]   = spc11_inst_done;//sparc 11
done[12]   = spc12_inst_done;//sparc 12
done[13]   = spc13_inst_done;//sparc 13
done[14]   = spc14_inst_done;//sparc 14
done[15]   = spc15_inst_done;//sparc 15
done[16]   = spc16_inst_done;//sparc 16
done[17]   = spc17_inst_done;//sparc 17
done[18]   = spc18_inst_done;//sparc 18
done[19]   = spc19_inst_done;//sparc 19
done[20]   = spc20_inst_done;//sparc 20
done[21]   = spc21_inst_done;//sparc 21
done[22]   = spc22_inst_done;//sparc 22
done[23]   = spc23_inst_done;//sparc 23
done[24]   = spc24_inst_done;//sparc 24
done[25]   = spc25_inst_done;//sparc 25
done[26]   = spc26_inst_done;//sparc 26
done[27]   = spc27_inst_done;//sparc 27
done[28]   = spc28_inst_done;//sparc 28
done[29]   = spc29_inst_done;//sparc 29
done[30]   = spc30_inst_done;//sparc 30
done[31]   = spc31_inst_done;//sparc 31
done[32]   = spc32_inst_done;//sparc 32
done[33]   = spc33_inst_done;//sparc 33
done[34]   = spc34_inst_done;//sparc 34
done[35]   = spc35_inst_done;//sparc 35
done[36]   = spc36_inst_done;//sparc 36
done[37]   = spc37_inst_done;//sparc 37
done[38]   = spc38_inst_done;//sparc 38
done[39]   = spc39_inst_done;//sparc 39
done[40]   = spc40_inst_done;//sparc 40
done[41]   = spc41_inst_done;//sparc 41
done[42]   = spc42_inst_done;//sparc 42
done[43]   = spc43_inst_done;//sparc 43
done[44]   = spc44_inst_done;//sparc 44
done[45]   = spc45_inst_done;//sparc 45
done[46]   = spc46_inst_done;//sparc 46
done[47]   = spc47_inst_done;//sparc 47
done[48]   = spc48_inst_done;//sparc 48
done[49]   = spc49_inst_done;//sparc 49
done[50]   = spc50_inst_done;//sparc 50
done[51]   = spc51_inst_done;//sparc 51
done[52]   = spc52_inst_done;//sparc 52
done[53]   = spc53_inst_done;//sparc 53
done[54]   = spc54_inst_done;//sparc 54
done[55]   = spc55_inst_done;//sparc 55
done[56]   = spc56_inst_done;//sparc 56
done[57]   = spc57_inst_done;//sparc 57
done[58]   = spc58_inst_done;//sparc 58
done[59]   = spc59_inst_done;//sparc 59
done[60]   = spc60_inst_done;//sparc 60
done[61]   = spc61_inst_done;//sparc 61
done[62]   = spc62_inst_done;//sparc 62
done[63]   = spc63_inst_done;//sparc 63
done[64]   = spc64_inst_done;//sparc 64
done[65]   = spc65_inst_done;//sparc 65
done[66]   = spc66_inst_done;//sparc 66
done[67]   = spc67_inst_done;//sparc 67
done[68]   = spc68_inst_done;//sparc 68
done[69]   = spc69_inst_done;//sparc 69
done[70]   = spc70_inst_done;//sparc 70
done[71]   = spc71_inst_done;//sparc 71
done[72]   = spc72_inst_done;//sparc 72
done[73]   = spc73_inst_done;//sparc 73
done[74]   = spc74_inst_done;//sparc 74
done[75]   = spc75_inst_done;//sparc 75
done[76]   = spc76_inst_done;//sparc 76
done[77]   = spc77_inst_done;//sparc 77
done[78]   = spc78_inst_done;//sparc 78
done[79]   = spc79_inst_done;//sparc 79
done[80]   = spc80_inst_done;//sparc 80
done[81]   = spc81_inst_done;//sparc 81
done[82]   = spc82_inst_done;//sparc 82
done[83]   = spc83_inst_done;//sparc 83
done[84]   = spc84_inst_done;//sparc 84
done[85]   = spc85_inst_done;//sparc 85
done[86]   = spc86_inst_done;//sparc 86
done[87]   = spc87_inst_done;//sparc 87
done[88]   = spc88_inst_done;//sparc 88
done[89]   = spc89_inst_done;//sparc 89
done[90]   = spc90_inst_done;//sparc 90
done[91]   = spc91_inst_done;//sparc 91
done[92]   = spc92_inst_done;//sparc 92
done[93]   = spc93_inst_done;//sparc 93
done[94]   = spc94_inst_done;//sparc 94
done[95]   = spc95_inst_done;//sparc 95
done[96]   = spc96_inst_done;//sparc 96
done[97]   = spc97_inst_done;//sparc 97
done[98]   = spc98_inst_done;//sparc 98
done[99]   = spc99_inst_done;//sparc 99
done[100]   = spc100_inst_done;//sparc 100
done[101]   = spc101_inst_done;//sparc 101
done[102]   = spc102_inst_done;//sparc 102
done[103]   = spc103_inst_done;//sparc 103
done[104]   = spc104_inst_done;//sparc 104
done[105]   = spc105_inst_done;//sparc 105
done[106]   = spc106_inst_done;//sparc 106
done[107]   = spc107_inst_done;//sparc 107
done[108]   = spc108_inst_done;//sparc 108
done[109]   = spc109_inst_done;//sparc 109
done[110]   = spc110_inst_done;//sparc 110
done[111]   = spc111_inst_done;//sparc 111
done[112]   = spc112_inst_done;//sparc 112
done[113]   = spc113_inst_done;//sparc 113
done[114]   = spc114_inst_done;//sparc 114
done[115]   = spc115_inst_done;//sparc 115
done[116]   = spc116_inst_done;//sparc 116
done[117]   = spc117_inst_done;//sparc 117
done[118]   = spc118_inst_done;//sparc 118
done[119]   = spc119_inst_done;//sparc 119
done[120]   = spc120_inst_done;//sparc 120
done[121]   = spc121_inst_done;//sparc 121
done[122]   = spc122_inst_done;//sparc 122
done[123]   = spc123_inst_done;//sparc 123
done[124]   = spc124_inst_done;//sparc 124
done[125]   = spc125_inst_done;//sparc 125
done[126]   = spc126_inst_done;//sparc 126
done[127]   = spc127_inst_done;//sparc 127
done[128]   = spc128_inst_done;//sparc 128
done[129]   = spc129_inst_done;//sparc 129
done[130]   = spc130_inst_done;//sparc 130
done[131]   = spc131_inst_done;//sparc 131
done[132]   = spc132_inst_done;//sparc 132
done[133]   = spc133_inst_done;//sparc 133
done[134]   = spc134_inst_done;//sparc 134
done[135]   = spc135_inst_done;//sparc 135
done[136]   = spc136_inst_done;//sparc 136
done[137]   = spc137_inst_done;//sparc 137
done[138]   = spc138_inst_done;//sparc 138
done[139]   = spc139_inst_done;//sparc 139
done[140]   = spc140_inst_done;//sparc 140
done[141]   = spc141_inst_done;//sparc 141
done[142]   = spc142_inst_done;//sparc 142
done[143]   = spc143_inst_done;//sparc 143
done[144]   = spc144_inst_done;//sparc 144
done[145]   = spc145_inst_done;//sparc 145
done[146]   = spc146_inst_done;//sparc 146
done[147]   = spc147_inst_done;//sparc 147
done[148]   = spc148_inst_done;//sparc 148
done[149]   = spc149_inst_done;//sparc 149
done[150]   = spc150_inst_done;//sparc 150
done[151]   = spc151_inst_done;//sparc 151
done[152]   = spc152_inst_done;//sparc 152
done[153]   = spc153_inst_done;//sparc 153
done[154]   = spc154_inst_done;//sparc 154
done[155]   = spc155_inst_done;//sparc 155
done[156]   = spc156_inst_done;//sparc 156
done[157]   = spc157_inst_done;//sparc 157
done[158]   = spc158_inst_done;//sparc 158
done[159]   = spc159_inst_done;//sparc 159
done[160]   = spc160_inst_done;//sparc 160
done[161]   = spc161_inst_done;//sparc 161
done[162]   = spc162_inst_done;//sparc 162
done[163]   = spc163_inst_done;//sparc 163
done[164]   = spc164_inst_done;//sparc 164
done[165]   = spc165_inst_done;//sparc 165
done[166]   = spc166_inst_done;//sparc 166
done[167]   = spc167_inst_done;//sparc 167
done[168]   = spc168_inst_done;//sparc 168
done[169]   = spc169_inst_done;//sparc 169
done[170]   = spc170_inst_done;//sparc 170
done[171]   = spc171_inst_done;//sparc 171
done[172]   = spc172_inst_done;//sparc 172
done[173]   = spc173_inst_done;//sparc 173
done[174]   = spc174_inst_done;//sparc 174
done[175]   = spc175_inst_done;//sparc 175
done[176]   = spc176_inst_done;//sparc 176
done[177]   = spc177_inst_done;//sparc 177
done[178]   = spc178_inst_done;//sparc 178
done[179]   = spc179_inst_done;//sparc 179
done[180]   = spc180_inst_done;//sparc 180
done[181]   = spc181_inst_done;//sparc 181
done[182]   = spc182_inst_done;//sparc 182
done[183]   = spc183_inst_done;//sparc 183
done[184]   = spc184_inst_done;//sparc 184
done[185]   = spc185_inst_done;//sparc 185
done[186]   = spc186_inst_done;//sparc 186
done[187]   = spc187_inst_done;//sparc 187
done[188]   = spc188_inst_done;//sparc 188
done[189]   = spc189_inst_done;//sparc 189
done[190]   = spc190_inst_done;//sparc 190
done[191]   = spc191_inst_done;//sparc 191
done[192]   = spc192_inst_done;//sparc 192
done[193]   = spc193_inst_done;//sparc 193
done[194]   = spc194_inst_done;//sparc 194
done[195]   = spc195_inst_done;//sparc 195
done[196]   = spc196_inst_done;//sparc 196
done[197]   = spc197_inst_done;//sparc 197
done[198]   = spc198_inst_done;//sparc 198
done[199]   = spc199_inst_done;//sparc 199
done[200]   = spc200_inst_done;//sparc 200
done[201]   = spc201_inst_done;//sparc 201
done[202]   = spc202_inst_done;//sparc 202
done[203]   = spc203_inst_done;//sparc 203
done[204]   = spc204_inst_done;//sparc 204
done[205]   = spc205_inst_done;//sparc 205
done[206]   = spc206_inst_done;//sparc 206
done[207]   = spc207_inst_done;//sparc 207
done[208]   = spc208_inst_done;//sparc 208
done[209]   = spc209_inst_done;//sparc 209
done[210]   = spc210_inst_done;//sparc 210
done[211]   = spc211_inst_done;//sparc 211
done[212]   = spc212_inst_done;//sparc 212
done[213]   = spc213_inst_done;//sparc 213
done[214]   = spc214_inst_done;//sparc 214
done[215]   = spc215_inst_done;//sparc 215
done[216]   = spc216_inst_done;//sparc 216
done[217]   = spc217_inst_done;//sparc 217
done[218]   = spc218_inst_done;//sparc 218
done[219]   = spc219_inst_done;//sparc 219
done[220]   = spc220_inst_done;//sparc 220
done[221]   = spc221_inst_done;//sparc 221
done[222]   = spc222_inst_done;//sparc 222
done[223]   = spc223_inst_done;//sparc 223
done[224]   = spc224_inst_done;//sparc 224
done[225]   = spc225_inst_done;//sparc 225
done[226]   = spc226_inst_done;//sparc 226
done[227]   = spc227_inst_done;//sparc 227
done[228]   = spc228_inst_done;//sparc 228
done[229]   = spc229_inst_done;//sparc 229
done[230]   = spc230_inst_done;//sparc 230
done[231]   = spc231_inst_done;//sparc 231
done[232]   = spc232_inst_done;//sparc 232
done[233]   = spc233_inst_done;//sparc 233
done[234]   = spc234_inst_done;//sparc 234
done[235]   = spc235_inst_done;//sparc 235
done[236]   = spc236_inst_done;//sparc 236
done[237]   = spc237_inst_done;//sparc 237
done[238]   = spc238_inst_done;//sparc 238
done[239]   = spc239_inst_done;//sparc 239
done[240]   = spc240_inst_done;//sparc 240
done[241]   = spc241_inst_done;//sparc 241
done[242]   = spc242_inst_done;//sparc 242
done[243]   = spc243_inst_done;//sparc 243
done[244]   = spc244_inst_done;//sparc 244
done[245]   = spc245_inst_done;//sparc 245
done[246]   = spc246_inst_done;//sparc 246
done[247]   = spc247_inst_done;//sparc 247
done[248]   = spc248_inst_done;//sparc 248
done[249]   = spc249_inst_done;//sparc 249
done[250]   = spc250_inst_done;//sparc 250
done[251]   = spc251_inst_done;//sparc 251
done[252]   = spc252_inst_done;//sparc 252
done[253]   = spc253_inst_done;//sparc 253
done[254]   = spc254_inst_done;//sparc 254
done[255]   = spc255_inst_done;//sparc 255
done[256]   = spc256_inst_done;//sparc 256
done[257]   = spc257_inst_done;//sparc 257
done[258]   = spc258_inst_done;//sparc 258
done[259]   = spc259_inst_done;//sparc 259
done[260]   = spc260_inst_done;//sparc 260
done[261]   = spc261_inst_done;//sparc 261
done[262]   = spc262_inst_done;//sparc 262
done[263]   = spc263_inst_done;//sparc 263
done[264]   = spc264_inst_done;//sparc 264
done[265]   = spc265_inst_done;//sparc 265
done[266]   = spc266_inst_done;//sparc 266
done[267]   = spc267_inst_done;//sparc 267
done[268]   = spc268_inst_done;//sparc 268
done[269]   = spc269_inst_done;//sparc 269
done[270]   = spc270_inst_done;//sparc 270
done[271]   = spc271_inst_done;//sparc 271
done[272]   = spc272_inst_done;//sparc 272
done[273]   = spc273_inst_done;//sparc 273
done[274]   = spc274_inst_done;//sparc 274
done[275]   = spc275_inst_done;//sparc 275
done[276]   = spc276_inst_done;//sparc 276
done[277]   = spc277_inst_done;//sparc 277
done[278]   = spc278_inst_done;//sparc 278
done[279]   = spc279_inst_done;//sparc 279
done[280]   = spc280_inst_done;//sparc 280
done[281]   = spc281_inst_done;//sparc 281
done[282]   = spc282_inst_done;//sparc 282
done[283]   = spc283_inst_done;//sparc 283
done[284]   = spc284_inst_done;//sparc 284
done[285]   = spc285_inst_done;//sparc 285
done[286]   = spc286_inst_done;//sparc 286
done[287]   = spc287_inst_done;//sparc 287
done[288]   = spc288_inst_done;//sparc 288
done[289]   = spc289_inst_done;//sparc 289
done[290]   = spc290_inst_done;//sparc 290
done[291]   = spc291_inst_done;//sparc 291
done[292]   = spc292_inst_done;//sparc 292
done[293]   = spc293_inst_done;//sparc 293
done[294]   = spc294_inst_done;//sparc 294
done[295]   = spc295_inst_done;//sparc 295
done[296]   = spc296_inst_done;//sparc 296
done[297]   = spc297_inst_done;//sparc 297
done[298]   = spc298_inst_done;//sparc 298
done[299]   = spc299_inst_done;//sparc 299
done[300]   = spc300_inst_done;//sparc 300
done[301]   = spc301_inst_done;//sparc 301
done[302]   = spc302_inst_done;//sparc 302
done[303]   = spc303_inst_done;//sparc 303
done[304]   = spc304_inst_done;//sparc 304
done[305]   = spc305_inst_done;//sparc 305
done[306]   = spc306_inst_done;//sparc 306
done[307]   = spc307_inst_done;//sparc 307
done[308]   = spc308_inst_done;//sparc 308
done[309]   = spc309_inst_done;//sparc 309
done[310]   = spc310_inst_done;//sparc 310
done[311]   = spc311_inst_done;//sparc 311
done[312]   = spc312_inst_done;//sparc 312
done[313]   = spc313_inst_done;//sparc 313
done[314]   = spc314_inst_done;//sparc 314
done[315]   = spc315_inst_done;//sparc 315
done[316]   = spc316_inst_done;//sparc 316
done[317]   = spc317_inst_done;//sparc 317
done[318]   = spc318_inst_done;//sparc 318
done[319]   = spc319_inst_done;//sparc 319
done[320]   = spc320_inst_done;//sparc 320
done[321]   = spc321_inst_done;//sparc 321
done[322]   = spc322_inst_done;//sparc 322
done[323]   = spc323_inst_done;//sparc 323
done[324]   = spc324_inst_done;//sparc 324
done[325]   = spc325_inst_done;//sparc 325
done[326]   = spc326_inst_done;//sparc 326
done[327]   = spc327_inst_done;//sparc 327
done[328]   = spc328_inst_done;//sparc 328
done[329]   = spc329_inst_done;//sparc 329
done[330]   = spc330_inst_done;//sparc 330
done[331]   = spc331_inst_done;//sparc 331
done[332]   = spc332_inst_done;//sparc 332
done[333]   = spc333_inst_done;//sparc 333
done[334]   = spc334_inst_done;//sparc 334
done[335]   = spc335_inst_done;//sparc 335
done[336]   = spc336_inst_done;//sparc 336
done[337]   = spc337_inst_done;//sparc 337
done[338]   = spc338_inst_done;//sparc 338
done[339]   = spc339_inst_done;//sparc 339
done[340]   = spc340_inst_done;//sparc 340
done[341]   = spc341_inst_done;//sparc 341
done[342]   = spc342_inst_done;//sparc 342
done[343]   = spc343_inst_done;//sparc 343
done[344]   = spc344_inst_done;//sparc 344
done[345]   = spc345_inst_done;//sparc 345
done[346]   = spc346_inst_done;//sparc 346
done[347]   = spc347_inst_done;//sparc 347
done[348]   = spc348_inst_done;//sparc 348
done[349]   = spc349_inst_done;//sparc 349
done[350]   = spc350_inst_done;//sparc 350
done[351]   = spc351_inst_done;//sparc 351
done[352]   = spc352_inst_done;//sparc 352
done[353]   = spc353_inst_done;//sparc 353
done[354]   = spc354_inst_done;//sparc 354
done[355]   = spc355_inst_done;//sparc 355
done[356]   = spc356_inst_done;//sparc 356
done[357]   = spc357_inst_done;//sparc 357
done[358]   = spc358_inst_done;//sparc 358
done[359]   = spc359_inst_done;//sparc 359
done[360]   = spc360_inst_done;//sparc 360
done[361]   = spc361_inst_done;//sparc 361
done[362]   = spc362_inst_done;//sparc 362
done[363]   = spc363_inst_done;//sparc 363
done[364]   = spc364_inst_done;//sparc 364
done[365]   = spc365_inst_done;//sparc 365
done[366]   = spc366_inst_done;//sparc 366
done[367]   = spc367_inst_done;//sparc 367
done[368]   = spc368_inst_done;//sparc 368
done[369]   = spc369_inst_done;//sparc 369
done[370]   = spc370_inst_done;//sparc 370
done[371]   = spc371_inst_done;//sparc 371
done[372]   = spc372_inst_done;//sparc 372
done[373]   = spc373_inst_done;//sparc 373
done[374]   = spc374_inst_done;//sparc 374
done[375]   = spc375_inst_done;//sparc 375
done[376]   = spc376_inst_done;//sparc 376
done[377]   = spc377_inst_done;//sparc 377
done[378]   = spc378_inst_done;//sparc 378
done[379]   = spc379_inst_done;//sparc 379
done[380]   = spc380_inst_done;//sparc 380
done[381]   = spc381_inst_done;//sparc 381
done[382]   = spc382_inst_done;//sparc 382
done[383]   = spc383_inst_done;//sparc 383
done[384]   = spc384_inst_done;//sparc 384
done[385]   = spc385_inst_done;//sparc 385
done[386]   = spc386_inst_done;//sparc 386
done[387]   = spc387_inst_done;//sparc 387
done[388]   = spc388_inst_done;//sparc 388
done[389]   = spc389_inst_done;//sparc 389
done[390]   = spc390_inst_done;//sparc 390
done[391]   = spc391_inst_done;//sparc 391
done[392]   = spc392_inst_done;//sparc 392
done[393]   = spc393_inst_done;//sparc 393
done[394]   = spc394_inst_done;//sparc 394
done[395]   = spc395_inst_done;//sparc 395
done[396]   = spc396_inst_done;//sparc 396
done[397]   = spc397_inst_done;//sparc 397
done[398]   = spc398_inst_done;//sparc 398
done[399]   = spc399_inst_done;//sparc 399
done[400]   = spc400_inst_done;//sparc 400
done[401]   = spc401_inst_done;//sparc 401
done[402]   = spc402_inst_done;//sparc 402
done[403]   = spc403_inst_done;//sparc 403
done[404]   = spc404_inst_done;//sparc 404
done[405]   = spc405_inst_done;//sparc 405
done[406]   = spc406_inst_done;//sparc 406
done[407]   = spc407_inst_done;//sparc 407
done[408]   = spc408_inst_done;//sparc 408
done[409]   = spc409_inst_done;//sparc 409
done[410]   = spc410_inst_done;//sparc 410
done[411]   = spc411_inst_done;//sparc 411
done[412]   = spc412_inst_done;//sparc 412
done[413]   = spc413_inst_done;//sparc 413
done[414]   = spc414_inst_done;//sparc 414
done[415]   = spc415_inst_done;//sparc 415
done[416]   = spc416_inst_done;//sparc 416
done[417]   = spc417_inst_done;//sparc 417
done[418]   = spc418_inst_done;//sparc 418
done[419]   = spc419_inst_done;//sparc 419
done[420]   = spc420_inst_done;//sparc 420
done[421]   = spc421_inst_done;//sparc 421
done[422]   = spc422_inst_done;//sparc 422
done[423]   = spc423_inst_done;//sparc 423
done[424]   = spc424_inst_done;//sparc 424
done[425]   = spc425_inst_done;//sparc 425
done[426]   = spc426_inst_done;//sparc 426
done[427]   = spc427_inst_done;//sparc 427
done[428]   = spc428_inst_done;//sparc 428
done[429]   = spc429_inst_done;//sparc 429
done[430]   = spc430_inst_done;//sparc 430
done[431]   = spc431_inst_done;//sparc 431
done[432]   = spc432_inst_done;//sparc 432
done[433]   = spc433_inst_done;//sparc 433
done[434]   = spc434_inst_done;//sparc 434
done[435]   = spc435_inst_done;//sparc 435
done[436]   = spc436_inst_done;//sparc 436
done[437]   = spc437_inst_done;//sparc 437
done[438]   = spc438_inst_done;//sparc 438
done[439]   = spc439_inst_done;//sparc 439
done[440]   = spc440_inst_done;//sparc 440
done[441]   = spc441_inst_done;//sparc 441
done[442]   = spc442_inst_done;//sparc 442
done[443]   = spc443_inst_done;//sparc 443
done[444]   = spc444_inst_done;//sparc 444
done[445]   = spc445_inst_done;//sparc 445
done[446]   = spc446_inst_done;//sparc 446
done[447]   = spc447_inst_done;//sparc 447
done[448]   = spc448_inst_done;//sparc 448
done[449]   = spc449_inst_done;//sparc 449
done[450]   = spc450_inst_done;//sparc 450
done[451]   = spc451_inst_done;//sparc 451
done[452]   = spc452_inst_done;//sparc 452
done[453]   = spc453_inst_done;//sparc 453
done[454]   = spc454_inst_done;//sparc 454
done[455]   = spc455_inst_done;//sparc 455
done[456]   = spc456_inst_done;//sparc 456
done[457]   = spc457_inst_done;//sparc 457
done[458]   = spc458_inst_done;//sparc 458
done[459]   = spc459_inst_done;//sparc 459
done[460]   = spc460_inst_done;//sparc 460
done[461]   = spc461_inst_done;//sparc 461
done[462]   = spc462_inst_done;//sparc 462
done[463]   = spc463_inst_done;//sparc 463
done[464]   = spc464_inst_done;//sparc 464
done[465]   = spc465_inst_done;//sparc 465
done[466]   = spc466_inst_done;//sparc 466
done[467]   = spc467_inst_done;//sparc 467
done[468]   = spc468_inst_done;//sparc 468
done[469]   = spc469_inst_done;//sparc 469
done[470]   = spc470_inst_done;//sparc 470
done[471]   = spc471_inst_done;//sparc 471
done[472]   = spc472_inst_done;//sparc 472
done[473]   = spc473_inst_done;//sparc 473
done[474]   = spc474_inst_done;//sparc 474
done[475]   = spc475_inst_done;//sparc 475
done[476]   = spc476_inst_done;//sparc 476
done[477]   = spc477_inst_done;//sparc 477
done[478]   = spc478_inst_done;//sparc 478
done[479]   = spc479_inst_done;//sparc 479
done[480]   = spc480_inst_done;//sparc 480
done[481]   = spc481_inst_done;//sparc 481
done[482]   = spc482_inst_done;//sparc 482
done[483]   = spc483_inst_done;//sparc 483
done[484]   = spc484_inst_done;//sparc 484
done[485]   = spc485_inst_done;//sparc 485
done[486]   = spc486_inst_done;//sparc 486
done[487]   = spc487_inst_done;//sparc 487
done[488]   = spc488_inst_done;//sparc 488
done[489]   = spc489_inst_done;//sparc 489
done[490]   = spc490_inst_done;//sparc 490
done[491]   = spc491_inst_done;//sparc 491
done[492]   = spc492_inst_done;//sparc 492
done[493]   = spc493_inst_done;//sparc 493
done[494]   = spc494_inst_done;//sparc 494
done[495]   = spc495_inst_done;//sparc 495
done[496]   = spc496_inst_done;//sparc 496
done[497]   = spc497_inst_done;//sparc 497
done[498]   = spc498_inst_done;//sparc 498
done[499]   = spc499_inst_done;//sparc 499
done[500]   = spc500_inst_done;//sparc 500
done[501]   = spc501_inst_done;//sparc 501
done[502]   = spc502_inst_done;//sparc 502
done[503]   = spc503_inst_done;//sparc 503
done[504]   = spc504_inst_done;//sparc 504
done[505]   = spc505_inst_done;//sparc 505
done[506]   = spc506_inst_done;//sparc 506
done[507]   = spc507_inst_done;//sparc 507
done[508]   = spc508_inst_done;//sparc 508
done[509]   = spc509_inst_done;//sparc 509
done[510]   = spc510_inst_done;//sparc 510
done[511]   = spc511_inst_done;//sparc 511
done[512]   = spc512_inst_done;//sparc 512
done[513]   = spc513_inst_done;//sparc 513
done[514]   = spc514_inst_done;//sparc 514
done[515]   = spc515_inst_done;//sparc 515
done[516]   = spc516_inst_done;//sparc 516
done[517]   = spc517_inst_done;//sparc 517
done[518]   = spc518_inst_done;//sparc 518
done[519]   = spc519_inst_done;//sparc 519
done[520]   = spc520_inst_done;//sparc 520
done[521]   = spc521_inst_done;//sparc 521
done[522]   = spc522_inst_done;//sparc 522
done[523]   = spc523_inst_done;//sparc 523
done[524]   = spc524_inst_done;//sparc 524
done[525]   = spc525_inst_done;//sparc 525
done[526]   = spc526_inst_done;//sparc 526
done[527]   = spc527_inst_done;//sparc 527
done[528]   = spc528_inst_done;//sparc 528
done[529]   = spc529_inst_done;//sparc 529
done[530]   = spc530_inst_done;//sparc 530
done[531]   = spc531_inst_done;//sparc 531
done[532]   = spc532_inst_done;//sparc 532
done[533]   = spc533_inst_done;//sparc 533
done[534]   = spc534_inst_done;//sparc 534
done[535]   = spc535_inst_done;//sparc 535
done[536]   = spc536_inst_done;//sparc 536
done[537]   = spc537_inst_done;//sparc 537
done[538]   = spc538_inst_done;//sparc 538
done[539]   = spc539_inst_done;//sparc 539
done[540]   = spc540_inst_done;//sparc 540
done[541]   = spc541_inst_done;//sparc 541
done[542]   = spc542_inst_done;//sparc 542
done[543]   = spc543_inst_done;//sparc 543
done[544]   = spc544_inst_done;//sparc 544
done[545]   = spc545_inst_done;//sparc 545
done[546]   = spc546_inst_done;//sparc 546
done[547]   = spc547_inst_done;//sparc 547
done[548]   = spc548_inst_done;//sparc 548
done[549]   = spc549_inst_done;//sparc 549
done[550]   = spc550_inst_done;//sparc 550
done[551]   = spc551_inst_done;//sparc 551
done[552]   = spc552_inst_done;//sparc 552
done[553]   = spc553_inst_done;//sparc 553
done[554]   = spc554_inst_done;//sparc 554
done[555]   = spc555_inst_done;//sparc 555
done[556]   = spc556_inst_done;//sparc 556
done[557]   = spc557_inst_done;//sparc 557
done[558]   = spc558_inst_done;//sparc 558
done[559]   = spc559_inst_done;//sparc 559
done[560]   = spc560_inst_done;//sparc 560
done[561]   = spc561_inst_done;//sparc 561
done[562]   = spc562_inst_done;//sparc 562
done[563]   = spc563_inst_done;//sparc 563
done[564]   = spc564_inst_done;//sparc 564
done[565]   = spc565_inst_done;//sparc 565
done[566]   = spc566_inst_done;//sparc 566
done[567]   = spc567_inst_done;//sparc 567
done[568]   = spc568_inst_done;//sparc 568
done[569]   = spc569_inst_done;//sparc 569
done[570]   = spc570_inst_done;//sparc 570
done[571]   = spc571_inst_done;//sparc 571
done[572]   = spc572_inst_done;//sparc 572
done[573]   = spc573_inst_done;//sparc 573
done[574]   = spc574_inst_done;//sparc 574
done[575]   = spc575_inst_done;//sparc 575
done[576]   = spc576_inst_done;//sparc 576
done[577]   = spc577_inst_done;//sparc 577
done[578]   = spc578_inst_done;//sparc 578
done[579]   = spc579_inst_done;//sparc 579
done[580]   = spc580_inst_done;//sparc 580
done[581]   = spc581_inst_done;//sparc 581
done[582]   = spc582_inst_done;//sparc 582
done[583]   = spc583_inst_done;//sparc 583
done[584]   = spc584_inst_done;//sparc 584
done[585]   = spc585_inst_done;//sparc 585
done[586]   = spc586_inst_done;//sparc 586
done[587]   = spc587_inst_done;//sparc 587
done[588]   = spc588_inst_done;//sparc 588
done[589]   = spc589_inst_done;//sparc 589
done[590]   = spc590_inst_done;//sparc 590
done[591]   = spc591_inst_done;//sparc 591
done[592]   = spc592_inst_done;//sparc 592
done[593]   = spc593_inst_done;//sparc 593
done[594]   = spc594_inst_done;//sparc 594
done[595]   = spc595_inst_done;//sparc 595
done[596]   = spc596_inst_done;//sparc 596
done[597]   = spc597_inst_done;//sparc 597
done[598]   = spc598_inst_done;//sparc 598
done[599]   = spc599_inst_done;//sparc 599
done[600]   = spc600_inst_done;//sparc 600
done[601]   = spc601_inst_done;//sparc 601
done[602]   = spc602_inst_done;//sparc 602
done[603]   = spc603_inst_done;//sparc 603
done[604]   = spc604_inst_done;//sparc 604
done[605]   = spc605_inst_done;//sparc 605
done[606]   = spc606_inst_done;//sparc 606
done[607]   = spc607_inst_done;//sparc 607
done[608]   = spc608_inst_done;//sparc 608
done[609]   = spc609_inst_done;//sparc 609
done[610]   = spc610_inst_done;//sparc 610
done[611]   = spc611_inst_done;//sparc 611
done[612]   = spc612_inst_done;//sparc 612
done[613]   = spc613_inst_done;//sparc 613
done[614]   = spc614_inst_done;//sparc 614
done[615]   = spc615_inst_done;//sparc 615
done[616]   = spc616_inst_done;//sparc 616
done[617]   = spc617_inst_done;//sparc 617
done[618]   = spc618_inst_done;//sparc 618
done[619]   = spc619_inst_done;//sparc 619
done[620]   = spc620_inst_done;//sparc 620
done[621]   = spc621_inst_done;//sparc 621
done[622]   = spc622_inst_done;//sparc 622
done[623]   = spc623_inst_done;//sparc 623
done[624]   = spc624_inst_done;//sparc 624
done[625]   = spc625_inst_done;//sparc 625
done[626]   = spc626_inst_done;//sparc 626
done[627]   = spc627_inst_done;//sparc 627
done[628]   = spc628_inst_done;//sparc 628
done[629]   = spc629_inst_done;//sparc 629
done[630]   = spc630_inst_done;//sparc 630
done[631]   = spc631_inst_done;//sparc 631
done[632]   = spc632_inst_done;//sparc 632
done[633]   = spc633_inst_done;//sparc 633
done[634]   = spc634_inst_done;//sparc 634
done[635]   = spc635_inst_done;//sparc 635
done[636]   = spc636_inst_done;//sparc 636
done[637]   = spc637_inst_done;//sparc 637
done[638]   = spc638_inst_done;//sparc 638
done[639]   = spc639_inst_done;//sparc 639
done[640]   = spc640_inst_done;//sparc 640
done[641]   = spc641_inst_done;//sparc 641
done[642]   = spc642_inst_done;//sparc 642
done[643]   = spc643_inst_done;//sparc 643
done[644]   = spc644_inst_done;//sparc 644
done[645]   = spc645_inst_done;//sparc 645
done[646]   = spc646_inst_done;//sparc 646
done[647]   = spc647_inst_done;//sparc 647
done[648]   = spc648_inst_done;//sparc 648
done[649]   = spc649_inst_done;//sparc 649
done[650]   = spc650_inst_done;//sparc 650
done[651]   = spc651_inst_done;//sparc 651
done[652]   = spc652_inst_done;//sparc 652
done[653]   = spc653_inst_done;//sparc 653
done[654]   = spc654_inst_done;//sparc 654
done[655]   = spc655_inst_done;//sparc 655
done[656]   = spc656_inst_done;//sparc 656
done[657]   = spc657_inst_done;//sparc 657
done[658]   = spc658_inst_done;//sparc 658
done[659]   = spc659_inst_done;//sparc 659
done[660]   = spc660_inst_done;//sparc 660
done[661]   = spc661_inst_done;//sparc 661
done[662]   = spc662_inst_done;//sparc 662
done[663]   = spc663_inst_done;//sparc 663
done[664]   = spc664_inst_done;//sparc 664
done[665]   = spc665_inst_done;//sparc 665
done[666]   = spc666_inst_done;//sparc 666
done[667]   = spc667_inst_done;//sparc 667
done[668]   = spc668_inst_done;//sparc 668
done[669]   = spc669_inst_done;//sparc 669
done[670]   = spc670_inst_done;//sparc 670
done[671]   = spc671_inst_done;//sparc 671
done[672]   = spc672_inst_done;//sparc 672
done[673]   = spc673_inst_done;//sparc 673
done[674]   = spc674_inst_done;//sparc 674
done[675]   = spc675_inst_done;//sparc 675
done[676]   = spc676_inst_done;//sparc 676
done[677]   = spc677_inst_done;//sparc 677
done[678]   = spc678_inst_done;//sparc 678
done[679]   = spc679_inst_done;//sparc 679
done[680]   = spc680_inst_done;//sparc 680
done[681]   = spc681_inst_done;//sparc 681
done[682]   = spc682_inst_done;//sparc 682
done[683]   = spc683_inst_done;//sparc 683
done[684]   = spc684_inst_done;//sparc 684
done[685]   = spc685_inst_done;//sparc 685
done[686]   = spc686_inst_done;//sparc 686
done[687]   = spc687_inst_done;//sparc 687
done[688]   = spc688_inst_done;//sparc 688
done[689]   = spc689_inst_done;//sparc 689
done[690]   = spc690_inst_done;//sparc 690
done[691]   = spc691_inst_done;//sparc 691
done[692]   = spc692_inst_done;//sparc 692
done[693]   = spc693_inst_done;//sparc 693
done[694]   = spc694_inst_done;//sparc 694
done[695]   = spc695_inst_done;//sparc 695
done[696]   = spc696_inst_done;//sparc 696
done[697]   = spc697_inst_done;//sparc 697
done[698]   = spc698_inst_done;//sparc 698
done[699]   = spc699_inst_done;//sparc 699
done[700]   = spc700_inst_done;//sparc 700
done[701]   = spc701_inst_done;//sparc 701
done[702]   = spc702_inst_done;//sparc 702
done[703]   = spc703_inst_done;//sparc 703
done[704]   = spc704_inst_done;//sparc 704
done[705]   = spc705_inst_done;//sparc 705
done[706]   = spc706_inst_done;//sparc 706
done[707]   = spc707_inst_done;//sparc 707
done[708]   = spc708_inst_done;//sparc 708
done[709]   = spc709_inst_done;//sparc 709
done[710]   = spc710_inst_done;//sparc 710
done[711]   = spc711_inst_done;//sparc 711
done[712]   = spc712_inst_done;//sparc 712
done[713]   = spc713_inst_done;//sparc 713
done[714]   = spc714_inst_done;//sparc 714
done[715]   = spc715_inst_done;//sparc 715
done[716]   = spc716_inst_done;//sparc 716
done[717]   = spc717_inst_done;//sparc 717
done[718]   = spc718_inst_done;//sparc 718
done[719]   = spc719_inst_done;//sparc 719
done[720]   = spc720_inst_done;//sparc 720
done[721]   = spc721_inst_done;//sparc 721
done[722]   = spc722_inst_done;//sparc 722
done[723]   = spc723_inst_done;//sparc 723
done[724]   = spc724_inst_done;//sparc 724
done[725]   = spc725_inst_done;//sparc 725
done[726]   = spc726_inst_done;//sparc 726
done[727]   = spc727_inst_done;//sparc 727
done[728]   = spc728_inst_done;//sparc 728
done[729]   = spc729_inst_done;//sparc 729
done[730]   = spc730_inst_done;//sparc 730
done[731]   = spc731_inst_done;//sparc 731
done[732]   = spc732_inst_done;//sparc 732
done[733]   = spc733_inst_done;//sparc 733
done[734]   = spc734_inst_done;//sparc 734
done[735]   = spc735_inst_done;//sparc 735
done[736]   = spc736_inst_done;//sparc 736
done[737]   = spc737_inst_done;//sparc 737
done[738]   = spc738_inst_done;//sparc 738
done[739]   = spc739_inst_done;//sparc 739
done[740]   = spc740_inst_done;//sparc 740
done[741]   = spc741_inst_done;//sparc 741
done[742]   = spc742_inst_done;//sparc 742
done[743]   = spc743_inst_done;//sparc 743
done[744]   = spc744_inst_done;//sparc 744
done[745]   = spc745_inst_done;//sparc 745
done[746]   = spc746_inst_done;//sparc 746
done[747]   = spc747_inst_done;//sparc 747
done[748]   = spc748_inst_done;//sparc 748
done[749]   = spc749_inst_done;//sparc 749
done[750]   = spc750_inst_done;//sparc 750
done[751]   = spc751_inst_done;//sparc 751
done[752]   = spc752_inst_done;//sparc 752
done[753]   = spc753_inst_done;//sparc 753
done[754]   = spc754_inst_done;//sparc 754
done[755]   = spc755_inst_done;//sparc 755
done[756]   = spc756_inst_done;//sparc 756
done[757]   = spc757_inst_done;//sparc 757
done[758]   = spc758_inst_done;//sparc 758
done[759]   = spc759_inst_done;//sparc 759
done[760]   = spc760_inst_done;//sparc 760
done[761]   = spc761_inst_done;//sparc 761
done[762]   = spc762_inst_done;//sparc 762
done[763]   = spc763_inst_done;//sparc 763
done[764]   = spc764_inst_done;//sparc 764
done[765]   = spc765_inst_done;//sparc 765
done[766]   = spc766_inst_done;//sparc 766
done[767]   = spc767_inst_done;//sparc 767
done[768]   = spc768_inst_done;//sparc 768
done[769]   = spc769_inst_done;//sparc 769
done[770]   = spc770_inst_done;//sparc 770
done[771]   = spc771_inst_done;//sparc 771
done[772]   = spc772_inst_done;//sparc 772
done[773]   = spc773_inst_done;//sparc 773
done[774]   = spc774_inst_done;//sparc 774
done[775]   = spc775_inst_done;//sparc 775
done[776]   = spc776_inst_done;//sparc 776
done[777]   = spc777_inst_done;//sparc 777
done[778]   = spc778_inst_done;//sparc 778
done[779]   = spc779_inst_done;//sparc 779
done[780]   = spc780_inst_done;//sparc 780
done[781]   = spc781_inst_done;//sparc 781
done[782]   = spc782_inst_done;//sparc 782
done[783]   = spc783_inst_done;//sparc 783
done[784]   = spc784_inst_done;//sparc 784
done[785]   = spc785_inst_done;//sparc 785
done[786]   = spc786_inst_done;//sparc 786
done[787]   = spc787_inst_done;//sparc 787
done[788]   = spc788_inst_done;//sparc 788
done[789]   = spc789_inst_done;//sparc 789
done[790]   = spc790_inst_done;//sparc 790
done[791]   = spc791_inst_done;//sparc 791
done[792]   = spc792_inst_done;//sparc 792
done[793]   = spc793_inst_done;//sparc 793
done[794]   = spc794_inst_done;//sparc 794
done[795]   = spc795_inst_done;//sparc 795
done[796]   = spc796_inst_done;//sparc 796
done[797]   = spc797_inst_done;//sparc 797
done[798]   = spc798_inst_done;//sparc 798
done[799]   = spc799_inst_done;//sparc 799
done[800]   = spc800_inst_done;//sparc 800
done[801]   = spc801_inst_done;//sparc 801
done[802]   = spc802_inst_done;//sparc 802
done[803]   = spc803_inst_done;//sparc 803
done[804]   = spc804_inst_done;//sparc 804
done[805]   = spc805_inst_done;//sparc 805
done[806]   = spc806_inst_done;//sparc 806
done[807]   = spc807_inst_done;//sparc 807
done[808]   = spc808_inst_done;//sparc 808
done[809]   = spc809_inst_done;//sparc 809
done[810]   = spc810_inst_done;//sparc 810
done[811]   = spc811_inst_done;//sparc 811
done[812]   = spc812_inst_done;//sparc 812
done[813]   = spc813_inst_done;//sparc 813
done[814]   = spc814_inst_done;//sparc 814
done[815]   = spc815_inst_done;//sparc 815
done[816]   = spc816_inst_done;//sparc 816
done[817]   = spc817_inst_done;//sparc 817
done[818]   = spc818_inst_done;//sparc 818
done[819]   = spc819_inst_done;//sparc 819
done[820]   = spc820_inst_done;//sparc 820
done[821]   = spc821_inst_done;//sparc 821
done[822]   = spc822_inst_done;//sparc 822
done[823]   = spc823_inst_done;//sparc 823
done[824]   = spc824_inst_done;//sparc 824
done[825]   = spc825_inst_done;//sparc 825
done[826]   = spc826_inst_done;//sparc 826
done[827]   = spc827_inst_done;//sparc 827
done[828]   = spc828_inst_done;//sparc 828
done[829]   = spc829_inst_done;//sparc 829
done[830]   = spc830_inst_done;//sparc 830
done[831]   = spc831_inst_done;//sparc 831
done[832]   = spc832_inst_done;//sparc 832
done[833]   = spc833_inst_done;//sparc 833
done[834]   = spc834_inst_done;//sparc 834
done[835]   = spc835_inst_done;//sparc 835
done[836]   = spc836_inst_done;//sparc 836
done[837]   = spc837_inst_done;//sparc 837
done[838]   = spc838_inst_done;//sparc 838
done[839]   = spc839_inst_done;//sparc 839
done[840]   = spc840_inst_done;//sparc 840
done[841]   = spc841_inst_done;//sparc 841
done[842]   = spc842_inst_done;//sparc 842
done[843]   = spc843_inst_done;//sparc 843
done[844]   = spc844_inst_done;//sparc 844
done[845]   = spc845_inst_done;//sparc 845
done[846]   = spc846_inst_done;//sparc 846
done[847]   = spc847_inst_done;//sparc 847
done[848]   = spc848_inst_done;//sparc 848
done[849]   = spc849_inst_done;//sparc 849
done[850]   = spc850_inst_done;//sparc 850
done[851]   = spc851_inst_done;//sparc 851
done[852]   = spc852_inst_done;//sparc 852
done[853]   = spc853_inst_done;//sparc 853
done[854]   = spc854_inst_done;//sparc 854
done[855]   = spc855_inst_done;//sparc 855
done[856]   = spc856_inst_done;//sparc 856
done[857]   = spc857_inst_done;//sparc 857
done[858]   = spc858_inst_done;//sparc 858
done[859]   = spc859_inst_done;//sparc 859
done[860]   = spc860_inst_done;//sparc 860
done[861]   = spc861_inst_done;//sparc 861
done[862]   = spc862_inst_done;//sparc 862
done[863]   = spc863_inst_done;//sparc 863
done[864]   = spc864_inst_done;//sparc 864
done[865]   = spc865_inst_done;//sparc 865
done[866]   = spc866_inst_done;//sparc 866
done[867]   = spc867_inst_done;//sparc 867
done[868]   = spc868_inst_done;//sparc 868
done[869]   = spc869_inst_done;//sparc 869
done[870]   = spc870_inst_done;//sparc 870
done[871]   = spc871_inst_done;//sparc 871
done[872]   = spc872_inst_done;//sparc 872
done[873]   = spc873_inst_done;//sparc 873
done[874]   = spc874_inst_done;//sparc 874
done[875]   = spc875_inst_done;//sparc 875
done[876]   = spc876_inst_done;//sparc 876
done[877]   = spc877_inst_done;//sparc 877
done[878]   = spc878_inst_done;//sparc 878
done[879]   = spc879_inst_done;//sparc 879
done[880]   = spc880_inst_done;//sparc 880
done[881]   = spc881_inst_done;//sparc 881
done[882]   = spc882_inst_done;//sparc 882
done[883]   = spc883_inst_done;//sparc 883
done[884]   = spc884_inst_done;//sparc 884
done[885]   = spc885_inst_done;//sparc 885
done[886]   = spc886_inst_done;//sparc 886
done[887]   = spc887_inst_done;//sparc 887
done[888]   = spc888_inst_done;//sparc 888
done[889]   = spc889_inst_done;//sparc 889
done[890]   = spc890_inst_done;//sparc 890
done[891]   = spc891_inst_done;//sparc 891
done[892]   = spc892_inst_done;//sparc 892
done[893]   = spc893_inst_done;//sparc 893
done[894]   = spc894_inst_done;//sparc 894
done[895]   = spc895_inst_done;//sparc 895
done[896]   = spc896_inst_done;//sparc 896
done[897]   = spc897_inst_done;//sparc 897
done[898]   = spc898_inst_done;//sparc 898
done[899]   = spc899_inst_done;//sparc 899
done[900]   = spc900_inst_done;//sparc 900
done[901]   = spc901_inst_done;//sparc 901
done[902]   = spc902_inst_done;//sparc 902
done[903]   = spc903_inst_done;//sparc 903
done[904]   = spc904_inst_done;//sparc 904
done[905]   = spc905_inst_done;//sparc 905
done[906]   = spc906_inst_done;//sparc 906
done[907]   = spc907_inst_done;//sparc 907
done[908]   = spc908_inst_done;//sparc 908
done[909]   = spc909_inst_done;//sparc 909
done[910]   = spc910_inst_done;//sparc 910
done[911]   = spc911_inst_done;//sparc 911
done[912]   = spc912_inst_done;//sparc 912
done[913]   = spc913_inst_done;//sparc 913
done[914]   = spc914_inst_done;//sparc 914
done[915]   = spc915_inst_done;//sparc 915
done[916]   = spc916_inst_done;//sparc 916
done[917]   = spc917_inst_done;//sparc 917
done[918]   = spc918_inst_done;//sparc 918
done[919]   = spc919_inst_done;//sparc 919
done[920]   = spc920_inst_done;//sparc 920
done[921]   = spc921_inst_done;//sparc 921
done[922]   = spc922_inst_done;//sparc 922
done[923]   = spc923_inst_done;//sparc 923
done[924]   = spc924_inst_done;//sparc 924
done[925]   = spc925_inst_done;//sparc 925
done[926]   = spc926_inst_done;//sparc 926
done[927]   = spc927_inst_done;//sparc 927
done[928]   = spc928_inst_done;//sparc 928
done[929]   = spc929_inst_done;//sparc 929
done[930]   = spc930_inst_done;//sparc 930
done[931]   = spc931_inst_done;//sparc 931
done[932]   = spc932_inst_done;//sparc 932
done[933]   = spc933_inst_done;//sparc 933
done[934]   = spc934_inst_done;//sparc 934
done[935]   = spc935_inst_done;//sparc 935
done[936]   = spc936_inst_done;//sparc 936
done[937]   = spc937_inst_done;//sparc 937
done[938]   = spc938_inst_done;//sparc 938
done[939]   = spc939_inst_done;//sparc 939
done[940]   = spc940_inst_done;//sparc 940
done[941]   = spc941_inst_done;//sparc 941
done[942]   = spc942_inst_done;//sparc 942
done[943]   = spc943_inst_done;//sparc 943
done[944]   = spc944_inst_done;//sparc 944
done[945]   = spc945_inst_done;//sparc 945
done[946]   = spc946_inst_done;//sparc 946
done[947]   = spc947_inst_done;//sparc 947
done[948]   = spc948_inst_done;//sparc 948
done[949]   = spc949_inst_done;//sparc 949
done[950]   = spc950_inst_done;//sparc 950
done[951]   = spc951_inst_done;//sparc 951
done[952]   = spc952_inst_done;//sparc 952
done[953]   = spc953_inst_done;//sparc 953
done[954]   = spc954_inst_done;//sparc 954
done[955]   = spc955_inst_done;//sparc 955
done[956]   = spc956_inst_done;//sparc 956
done[957]   = spc957_inst_done;//sparc 957
done[958]   = spc958_inst_done;//sparc 958
done[959]   = spc959_inst_done;//sparc 959
done[960]   = spc960_inst_done;//sparc 960
done[961]   = spc961_inst_done;//sparc 961
done[962]   = spc962_inst_done;//sparc 962
done[963]   = spc963_inst_done;//sparc 963
done[964]   = spc964_inst_done;//sparc 964
done[965]   = spc965_inst_done;//sparc 965
done[966]   = spc966_inst_done;//sparc 966
done[967]   = spc967_inst_done;//sparc 967
done[968]   = spc968_inst_done;//sparc 968
done[969]   = spc969_inst_done;//sparc 969
done[970]   = spc970_inst_done;//sparc 970
done[971]   = spc971_inst_done;//sparc 971
done[972]   = spc972_inst_done;//sparc 972
done[973]   = spc973_inst_done;//sparc 973
done[974]   = spc974_inst_done;//sparc 974
done[975]   = spc975_inst_done;//sparc 975
done[976]   = spc976_inst_done;//sparc 976
done[977]   = spc977_inst_done;//sparc 977
done[978]   = spc978_inst_done;//sparc 978
done[979]   = spc979_inst_done;//sparc 979
done[980]   = spc980_inst_done;//sparc 980
done[981]   = spc981_inst_done;//sparc 981
done[982]   = spc982_inst_done;//sparc 982
done[983]   = spc983_inst_done;//sparc 983
done[984]   = spc984_inst_done;//sparc 984
done[985]   = spc985_inst_done;//sparc 985
done[986]   = spc986_inst_done;//sparc 986
done[987]   = spc987_inst_done;//sparc 987
done[988]   = spc988_inst_done;//sparc 988
done[989]   = spc989_inst_done;//sparc 989
done[990]   = spc990_inst_done;//sparc 990
done[991]   = spc991_inst_done;//sparc 991
done[992]   = spc992_inst_done;//sparc 992
done[993]   = spc993_inst_done;//sparc 993
done[994]   = spc994_inst_done;//sparc 994
done[995]   = spc995_inst_done;//sparc 995
done[996]   = spc996_inst_done;//sparc 996
done[997]   = spc997_inst_done;//sparc 997
done[998]   = spc998_inst_done;//sparc 998
done[999]   = spc999_inst_done;//sparc 999
done[1000]   = spc1000_inst_done;//sparc 1000
done[1001]   = spc1001_inst_done;//sparc 1001
done[1002]   = spc1002_inst_done;//sparc 1002
done[1003]   = spc1003_inst_done;//sparc 1003
done[1004]   = spc1004_inst_done;//sparc 1004
done[1005]   = spc1005_inst_done;//sparc 1005
done[1006]   = spc1006_inst_done;//sparc 1006
done[1007]   = spc1007_inst_done;//sparc 1007
done[1008]   = spc1008_inst_done;//sparc 1008
done[1009]   = spc1009_inst_done;//sparc 1009
done[1010]   = spc1010_inst_done;//sparc 1010
done[1011]   = spc1011_inst_done;//sparc 1011
done[1012]   = spc1012_inst_done;//sparc 1012
done[1013]   = spc1013_inst_done;//sparc 1013
done[1014]   = spc1014_inst_done;//sparc 1014
done[1015]   = spc1015_inst_done;//sparc 1015
done[1016]   = spc1016_inst_done;//sparc 1016
done[1017]   = spc1017_inst_done;//sparc 1017
done[1018]   = spc1018_inst_done;//sparc 1018
done[1019]   = spc1019_inst_done;//sparc 1019
done[1020]   = spc1020_inst_done;//sparc 1020
done[1021]   = spc1021_inst_done;//sparc 1021
done[1022]   = spc1022_inst_done;//sparc 1022
done[1023]   = spc1023_inst_done;//sparc 1023


end



string linebuf0 = "";
logic hitMadPrint0 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc0_inst_done && ((spc0_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint0 = 1;
       linebuf0 = {linebuf0, spc0_phy_pc_w[8:1]};
       if (spc0_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 0, linebuf0);
          linebuf0 = "";
       end
    end else begin
       hitMadPrint0 = 0;
    end
  end
end


string linebuf1 = "";
logic hitMadPrint1 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc1_inst_done && ((spc1_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint1 = 1;
       linebuf1 = {linebuf1, spc1_phy_pc_w[8:1]};
       if (spc1_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 1, linebuf1);
          linebuf1 = "";
       end
    end else begin
       hitMadPrint1 = 0;
    end
  end
end


string linebuf2 = "";
logic hitMadPrint2 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc2_inst_done && ((spc2_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint2 = 1;
       linebuf2 = {linebuf2, spc2_phy_pc_w[8:1]};
       if (spc2_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 2, linebuf2);
          linebuf2 = "";
       end
    end else begin
       hitMadPrint2 = 0;
    end
  end
end


string linebuf3 = "";
logic hitMadPrint3 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc3_inst_done && ((spc3_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint3 = 1;
       linebuf3 = {linebuf3, spc3_phy_pc_w[8:1]};
       if (spc3_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 3, linebuf3);
          linebuf3 = "";
       end
    end else begin
       hitMadPrint3 = 0;
    end
  end
end


string linebuf4 = "";
logic hitMadPrint4 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc4_inst_done && ((spc4_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint4 = 1;
       linebuf4 = {linebuf4, spc4_phy_pc_w[8:1]};
       if (spc4_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 4, linebuf4);
          linebuf4 = "";
       end
    end else begin
       hitMadPrint4 = 0;
    end
  end
end


string linebuf5 = "";
logic hitMadPrint5 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc5_inst_done && ((spc5_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint5 = 1;
       linebuf5 = {linebuf5, spc5_phy_pc_w[8:1]};
       if (spc5_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 5, linebuf5);
          linebuf5 = "";
       end
    end else begin
       hitMadPrint5 = 0;
    end
  end
end


string linebuf6 = "";
logic hitMadPrint6 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc6_inst_done && ((spc6_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint6 = 1;
       linebuf6 = {linebuf6, spc6_phy_pc_w[8:1]};
       if (spc6_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 6, linebuf6);
          linebuf6 = "";
       end
    end else begin
       hitMadPrint6 = 0;
    end
  end
end


string linebuf7 = "";
logic hitMadPrint7 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc7_inst_done && ((spc7_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint7 = 1;
       linebuf7 = {linebuf7, spc7_phy_pc_w[8:1]};
       if (spc7_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 7, linebuf7);
          linebuf7 = "";
       end
    end else begin
       hitMadPrint7 = 0;
    end
  end
end


string linebuf8 = "";
logic hitMadPrint8 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc8_inst_done && ((spc8_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint8 = 1;
       linebuf8 = {linebuf8, spc8_phy_pc_w[8:1]};
       if (spc8_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 8, linebuf8);
          linebuf8 = "";
       end
    end else begin
       hitMadPrint8 = 0;
    end
  end
end


string linebuf9 = "";
logic hitMadPrint9 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc9_inst_done && ((spc9_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint9 = 1;
       linebuf9 = {linebuf9, spc9_phy_pc_w[8:1]};
       if (spc9_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 9, linebuf9);
          linebuf9 = "";
       end
    end else begin
       hitMadPrint9 = 0;
    end
  end
end


string linebuf10 = "";
logic hitMadPrint10 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc10_inst_done && ((spc10_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint10 = 1;
       linebuf10 = {linebuf10, spc10_phy_pc_w[8:1]};
       if (spc10_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 10, linebuf10);
          linebuf10 = "";
       end
    end else begin
       hitMadPrint10 = 0;
    end
  end
end


string linebuf11 = "";
logic hitMadPrint11 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc11_inst_done && ((spc11_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint11 = 1;
       linebuf11 = {linebuf11, spc11_phy_pc_w[8:1]};
       if (spc11_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 11, linebuf11);
          linebuf11 = "";
       end
    end else begin
       hitMadPrint11 = 0;
    end
  end
end


string linebuf12 = "";
logic hitMadPrint12 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc12_inst_done && ((spc12_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint12 = 1;
       linebuf12 = {linebuf12, spc12_phy_pc_w[8:1]};
       if (spc12_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 12, linebuf12);
          linebuf12 = "";
       end
    end else begin
       hitMadPrint12 = 0;
    end
  end
end


string linebuf13 = "";
logic hitMadPrint13 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc13_inst_done && ((spc13_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint13 = 1;
       linebuf13 = {linebuf13, spc13_phy_pc_w[8:1]};
       if (spc13_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 13, linebuf13);
          linebuf13 = "";
       end
    end else begin
       hitMadPrint13 = 0;
    end
  end
end


string linebuf14 = "";
logic hitMadPrint14 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc14_inst_done && ((spc14_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint14 = 1;
       linebuf14 = {linebuf14, spc14_phy_pc_w[8:1]};
       if (spc14_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 14, linebuf14);
          linebuf14 = "";
       end
    end else begin
       hitMadPrint14 = 0;
    end
  end
end


string linebuf15 = "";
logic hitMadPrint15 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc15_inst_done && ((spc15_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint15 = 1;
       linebuf15 = {linebuf15, spc15_phy_pc_w[8:1]};
       if (spc15_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 15, linebuf15);
          linebuf15 = "";
       end
    end else begin
       hitMadPrint15 = 0;
    end
  end
end


string linebuf16 = "";
logic hitMadPrint16 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc16_inst_done && ((spc16_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint16 = 1;
       linebuf16 = {linebuf16, spc16_phy_pc_w[8:1]};
       if (spc16_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 16, linebuf16);
          linebuf16 = "";
       end
    end else begin
       hitMadPrint16 = 0;
    end
  end
end


string linebuf17 = "";
logic hitMadPrint17 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc17_inst_done && ((spc17_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint17 = 1;
       linebuf17 = {linebuf17, spc17_phy_pc_w[8:1]};
       if (spc17_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 17, linebuf17);
          linebuf17 = "";
       end
    end else begin
       hitMadPrint17 = 0;
    end
  end
end


string linebuf18 = "";
logic hitMadPrint18 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc18_inst_done && ((spc18_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint18 = 1;
       linebuf18 = {linebuf18, spc18_phy_pc_w[8:1]};
       if (spc18_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 18, linebuf18);
          linebuf18 = "";
       end
    end else begin
       hitMadPrint18 = 0;
    end
  end
end


string linebuf19 = "";
logic hitMadPrint19 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc19_inst_done && ((spc19_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint19 = 1;
       linebuf19 = {linebuf19, spc19_phy_pc_w[8:1]};
       if (spc19_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 19, linebuf19);
          linebuf19 = "";
       end
    end else begin
       hitMadPrint19 = 0;
    end
  end
end


string linebuf20 = "";
logic hitMadPrint20 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc20_inst_done && ((spc20_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint20 = 1;
       linebuf20 = {linebuf20, spc20_phy_pc_w[8:1]};
       if (spc20_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 20, linebuf20);
          linebuf20 = "";
       end
    end else begin
       hitMadPrint20 = 0;
    end
  end
end


string linebuf21 = "";
logic hitMadPrint21 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc21_inst_done && ((spc21_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint21 = 1;
       linebuf21 = {linebuf21, spc21_phy_pc_w[8:1]};
       if (spc21_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 21, linebuf21);
          linebuf21 = "";
       end
    end else begin
       hitMadPrint21 = 0;
    end
  end
end


string linebuf22 = "";
logic hitMadPrint22 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc22_inst_done && ((spc22_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint22 = 1;
       linebuf22 = {linebuf22, spc22_phy_pc_w[8:1]};
       if (spc22_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 22, linebuf22);
          linebuf22 = "";
       end
    end else begin
       hitMadPrint22 = 0;
    end
  end
end


string linebuf23 = "";
logic hitMadPrint23 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc23_inst_done && ((spc23_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint23 = 1;
       linebuf23 = {linebuf23, spc23_phy_pc_w[8:1]};
       if (spc23_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 23, linebuf23);
          linebuf23 = "";
       end
    end else begin
       hitMadPrint23 = 0;
    end
  end
end


string linebuf24 = "";
logic hitMadPrint24 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc24_inst_done && ((spc24_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint24 = 1;
       linebuf24 = {linebuf24, spc24_phy_pc_w[8:1]};
       if (spc24_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 24, linebuf24);
          linebuf24 = "";
       end
    end else begin
       hitMadPrint24 = 0;
    end
  end
end


string linebuf25 = "";
logic hitMadPrint25 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc25_inst_done && ((spc25_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint25 = 1;
       linebuf25 = {linebuf25, spc25_phy_pc_w[8:1]};
       if (spc25_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 25, linebuf25);
          linebuf25 = "";
       end
    end else begin
       hitMadPrint25 = 0;
    end
  end
end


string linebuf26 = "";
logic hitMadPrint26 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc26_inst_done && ((spc26_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint26 = 1;
       linebuf26 = {linebuf26, spc26_phy_pc_w[8:1]};
       if (spc26_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 26, linebuf26);
          linebuf26 = "";
       end
    end else begin
       hitMadPrint26 = 0;
    end
  end
end


string linebuf27 = "";
logic hitMadPrint27 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc27_inst_done && ((spc27_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint27 = 1;
       linebuf27 = {linebuf27, spc27_phy_pc_w[8:1]};
       if (spc27_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 27, linebuf27);
          linebuf27 = "";
       end
    end else begin
       hitMadPrint27 = 0;
    end
  end
end


string linebuf28 = "";
logic hitMadPrint28 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc28_inst_done && ((spc28_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint28 = 1;
       linebuf28 = {linebuf28, spc28_phy_pc_w[8:1]};
       if (spc28_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 28, linebuf28);
          linebuf28 = "";
       end
    end else begin
       hitMadPrint28 = 0;
    end
  end
end


string linebuf29 = "";
logic hitMadPrint29 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc29_inst_done && ((spc29_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint29 = 1;
       linebuf29 = {linebuf29, spc29_phy_pc_w[8:1]};
       if (spc29_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 29, linebuf29);
          linebuf29 = "";
       end
    end else begin
       hitMadPrint29 = 0;
    end
  end
end


string linebuf30 = "";
logic hitMadPrint30 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc30_inst_done && ((spc30_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint30 = 1;
       linebuf30 = {linebuf30, spc30_phy_pc_w[8:1]};
       if (spc30_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 30, linebuf30);
          linebuf30 = "";
       end
    end else begin
       hitMadPrint30 = 0;
    end
  end
end


string linebuf31 = "";
logic hitMadPrint31 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc31_inst_done && ((spc31_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint31 = 1;
       linebuf31 = {linebuf31, spc31_phy_pc_w[8:1]};
       if (spc31_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 31, linebuf31);
          linebuf31 = "";
       end
    end else begin
       hitMadPrint31 = 0;
    end
  end
end


string linebuf32 = "";
logic hitMadPrint32 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc32_inst_done && ((spc32_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint32 = 1;
       linebuf32 = {linebuf32, spc32_phy_pc_w[8:1]};
       if (spc32_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 32, linebuf32);
          linebuf32 = "";
       end
    end else begin
       hitMadPrint32 = 0;
    end
  end
end


string linebuf33 = "";
logic hitMadPrint33 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc33_inst_done && ((spc33_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint33 = 1;
       linebuf33 = {linebuf33, spc33_phy_pc_w[8:1]};
       if (spc33_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 33, linebuf33);
          linebuf33 = "";
       end
    end else begin
       hitMadPrint33 = 0;
    end
  end
end


string linebuf34 = "";
logic hitMadPrint34 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc34_inst_done && ((spc34_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint34 = 1;
       linebuf34 = {linebuf34, spc34_phy_pc_w[8:1]};
       if (spc34_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 34, linebuf34);
          linebuf34 = "";
       end
    end else begin
       hitMadPrint34 = 0;
    end
  end
end


string linebuf35 = "";
logic hitMadPrint35 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc35_inst_done && ((spc35_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint35 = 1;
       linebuf35 = {linebuf35, spc35_phy_pc_w[8:1]};
       if (spc35_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 35, linebuf35);
          linebuf35 = "";
       end
    end else begin
       hitMadPrint35 = 0;
    end
  end
end


string linebuf36 = "";
logic hitMadPrint36 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc36_inst_done && ((spc36_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint36 = 1;
       linebuf36 = {linebuf36, spc36_phy_pc_w[8:1]};
       if (spc36_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 36, linebuf36);
          linebuf36 = "";
       end
    end else begin
       hitMadPrint36 = 0;
    end
  end
end


string linebuf37 = "";
logic hitMadPrint37 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc37_inst_done && ((spc37_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint37 = 1;
       linebuf37 = {linebuf37, spc37_phy_pc_w[8:1]};
       if (spc37_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 37, linebuf37);
          linebuf37 = "";
       end
    end else begin
       hitMadPrint37 = 0;
    end
  end
end


string linebuf38 = "";
logic hitMadPrint38 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc38_inst_done && ((spc38_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint38 = 1;
       linebuf38 = {linebuf38, spc38_phy_pc_w[8:1]};
       if (spc38_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 38, linebuf38);
          linebuf38 = "";
       end
    end else begin
       hitMadPrint38 = 0;
    end
  end
end


string linebuf39 = "";
logic hitMadPrint39 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc39_inst_done && ((spc39_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint39 = 1;
       linebuf39 = {linebuf39, spc39_phy_pc_w[8:1]};
       if (spc39_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 39, linebuf39);
          linebuf39 = "";
       end
    end else begin
       hitMadPrint39 = 0;
    end
  end
end


string linebuf40 = "";
logic hitMadPrint40 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc40_inst_done && ((spc40_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint40 = 1;
       linebuf40 = {linebuf40, spc40_phy_pc_w[8:1]};
       if (spc40_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 40, linebuf40);
          linebuf40 = "";
       end
    end else begin
       hitMadPrint40 = 0;
    end
  end
end


string linebuf41 = "";
logic hitMadPrint41 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc41_inst_done && ((spc41_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint41 = 1;
       linebuf41 = {linebuf41, spc41_phy_pc_w[8:1]};
       if (spc41_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 41, linebuf41);
          linebuf41 = "";
       end
    end else begin
       hitMadPrint41 = 0;
    end
  end
end


string linebuf42 = "";
logic hitMadPrint42 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc42_inst_done && ((spc42_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint42 = 1;
       linebuf42 = {linebuf42, spc42_phy_pc_w[8:1]};
       if (spc42_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 42, linebuf42);
          linebuf42 = "";
       end
    end else begin
       hitMadPrint42 = 0;
    end
  end
end


string linebuf43 = "";
logic hitMadPrint43 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc43_inst_done && ((spc43_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint43 = 1;
       linebuf43 = {linebuf43, spc43_phy_pc_w[8:1]};
       if (spc43_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 43, linebuf43);
          linebuf43 = "";
       end
    end else begin
       hitMadPrint43 = 0;
    end
  end
end


string linebuf44 = "";
logic hitMadPrint44 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc44_inst_done && ((spc44_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint44 = 1;
       linebuf44 = {linebuf44, spc44_phy_pc_w[8:1]};
       if (spc44_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 44, linebuf44);
          linebuf44 = "";
       end
    end else begin
       hitMadPrint44 = 0;
    end
  end
end


string linebuf45 = "";
logic hitMadPrint45 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc45_inst_done && ((spc45_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint45 = 1;
       linebuf45 = {linebuf45, spc45_phy_pc_w[8:1]};
       if (spc45_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 45, linebuf45);
          linebuf45 = "";
       end
    end else begin
       hitMadPrint45 = 0;
    end
  end
end


string linebuf46 = "";
logic hitMadPrint46 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc46_inst_done && ((spc46_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint46 = 1;
       linebuf46 = {linebuf46, spc46_phy_pc_w[8:1]};
       if (spc46_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 46, linebuf46);
          linebuf46 = "";
       end
    end else begin
       hitMadPrint46 = 0;
    end
  end
end


string linebuf47 = "";
logic hitMadPrint47 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc47_inst_done && ((spc47_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint47 = 1;
       linebuf47 = {linebuf47, spc47_phy_pc_w[8:1]};
       if (spc47_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 47, linebuf47);
          linebuf47 = "";
       end
    end else begin
       hitMadPrint47 = 0;
    end
  end
end


string linebuf48 = "";
logic hitMadPrint48 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc48_inst_done && ((spc48_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint48 = 1;
       linebuf48 = {linebuf48, spc48_phy_pc_w[8:1]};
       if (spc48_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 48, linebuf48);
          linebuf48 = "";
       end
    end else begin
       hitMadPrint48 = 0;
    end
  end
end


string linebuf49 = "";
logic hitMadPrint49 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc49_inst_done && ((spc49_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint49 = 1;
       linebuf49 = {linebuf49, spc49_phy_pc_w[8:1]};
       if (spc49_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 49, linebuf49);
          linebuf49 = "";
       end
    end else begin
       hitMadPrint49 = 0;
    end
  end
end


string linebuf50 = "";
logic hitMadPrint50 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc50_inst_done && ((spc50_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint50 = 1;
       linebuf50 = {linebuf50, spc50_phy_pc_w[8:1]};
       if (spc50_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 50, linebuf50);
          linebuf50 = "";
       end
    end else begin
       hitMadPrint50 = 0;
    end
  end
end


string linebuf51 = "";
logic hitMadPrint51 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc51_inst_done && ((spc51_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint51 = 1;
       linebuf51 = {linebuf51, spc51_phy_pc_w[8:1]};
       if (spc51_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 51, linebuf51);
          linebuf51 = "";
       end
    end else begin
       hitMadPrint51 = 0;
    end
  end
end


string linebuf52 = "";
logic hitMadPrint52 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc52_inst_done && ((spc52_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint52 = 1;
       linebuf52 = {linebuf52, spc52_phy_pc_w[8:1]};
       if (spc52_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 52, linebuf52);
          linebuf52 = "";
       end
    end else begin
       hitMadPrint52 = 0;
    end
  end
end


string linebuf53 = "";
logic hitMadPrint53 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc53_inst_done && ((spc53_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint53 = 1;
       linebuf53 = {linebuf53, spc53_phy_pc_w[8:1]};
       if (spc53_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 53, linebuf53);
          linebuf53 = "";
       end
    end else begin
       hitMadPrint53 = 0;
    end
  end
end


string linebuf54 = "";
logic hitMadPrint54 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc54_inst_done && ((spc54_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint54 = 1;
       linebuf54 = {linebuf54, spc54_phy_pc_w[8:1]};
       if (spc54_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 54, linebuf54);
          linebuf54 = "";
       end
    end else begin
       hitMadPrint54 = 0;
    end
  end
end


string linebuf55 = "";
logic hitMadPrint55 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc55_inst_done && ((spc55_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint55 = 1;
       linebuf55 = {linebuf55, spc55_phy_pc_w[8:1]};
       if (spc55_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 55, linebuf55);
          linebuf55 = "";
       end
    end else begin
       hitMadPrint55 = 0;
    end
  end
end


string linebuf56 = "";
logic hitMadPrint56 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc56_inst_done && ((spc56_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint56 = 1;
       linebuf56 = {linebuf56, spc56_phy_pc_w[8:1]};
       if (spc56_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 56, linebuf56);
          linebuf56 = "";
       end
    end else begin
       hitMadPrint56 = 0;
    end
  end
end


string linebuf57 = "";
logic hitMadPrint57 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc57_inst_done && ((spc57_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint57 = 1;
       linebuf57 = {linebuf57, spc57_phy_pc_w[8:1]};
       if (spc57_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 57, linebuf57);
          linebuf57 = "";
       end
    end else begin
       hitMadPrint57 = 0;
    end
  end
end


string linebuf58 = "";
logic hitMadPrint58 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc58_inst_done && ((spc58_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint58 = 1;
       linebuf58 = {linebuf58, spc58_phy_pc_w[8:1]};
       if (spc58_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 58, linebuf58);
          linebuf58 = "";
       end
    end else begin
       hitMadPrint58 = 0;
    end
  end
end


string linebuf59 = "";
logic hitMadPrint59 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc59_inst_done && ((spc59_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint59 = 1;
       linebuf59 = {linebuf59, spc59_phy_pc_w[8:1]};
       if (spc59_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 59, linebuf59);
          linebuf59 = "";
       end
    end else begin
       hitMadPrint59 = 0;
    end
  end
end


string linebuf60 = "";
logic hitMadPrint60 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc60_inst_done && ((spc60_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint60 = 1;
       linebuf60 = {linebuf60, spc60_phy_pc_w[8:1]};
       if (spc60_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 60, linebuf60);
          linebuf60 = "";
       end
    end else begin
       hitMadPrint60 = 0;
    end
  end
end


string linebuf61 = "";
logic hitMadPrint61 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc61_inst_done && ((spc61_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint61 = 1;
       linebuf61 = {linebuf61, spc61_phy_pc_w[8:1]};
       if (spc61_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 61, linebuf61);
          linebuf61 = "";
       end
    end else begin
       hitMadPrint61 = 0;
    end
  end
end


string linebuf62 = "";
logic hitMadPrint62 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc62_inst_done && ((spc62_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint62 = 1;
       linebuf62 = {linebuf62, spc62_phy_pc_w[8:1]};
       if (spc62_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 62, linebuf62);
          linebuf62 = "";
       end
    end else begin
       hitMadPrint62 = 0;
    end
  end
end


string linebuf63 = "";
logic hitMadPrint63 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc63_inst_done && ((spc63_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint63 = 1;
       linebuf63 = {linebuf63, spc63_phy_pc_w[8:1]};
       if (spc63_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 63, linebuf63);
          linebuf63 = "";
       end
    end else begin
       hitMadPrint63 = 0;
    end
  end
end


string linebuf64 = "";
logic hitMadPrint64 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc64_inst_done && ((spc64_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint64 = 1;
       linebuf64 = {linebuf64, spc64_phy_pc_w[8:1]};
       if (spc64_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 64, linebuf64);
          linebuf64 = "";
       end
    end else begin
       hitMadPrint64 = 0;
    end
  end
end


string linebuf65 = "";
logic hitMadPrint65 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc65_inst_done && ((spc65_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint65 = 1;
       linebuf65 = {linebuf65, spc65_phy_pc_w[8:1]};
       if (spc65_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 65, linebuf65);
          linebuf65 = "";
       end
    end else begin
       hitMadPrint65 = 0;
    end
  end
end


string linebuf66 = "";
logic hitMadPrint66 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc66_inst_done && ((spc66_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint66 = 1;
       linebuf66 = {linebuf66, spc66_phy_pc_w[8:1]};
       if (spc66_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 66, linebuf66);
          linebuf66 = "";
       end
    end else begin
       hitMadPrint66 = 0;
    end
  end
end


string linebuf67 = "";
logic hitMadPrint67 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc67_inst_done && ((spc67_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint67 = 1;
       linebuf67 = {linebuf67, spc67_phy_pc_w[8:1]};
       if (spc67_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 67, linebuf67);
          linebuf67 = "";
       end
    end else begin
       hitMadPrint67 = 0;
    end
  end
end


string linebuf68 = "";
logic hitMadPrint68 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc68_inst_done && ((spc68_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint68 = 1;
       linebuf68 = {linebuf68, spc68_phy_pc_w[8:1]};
       if (spc68_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 68, linebuf68);
          linebuf68 = "";
       end
    end else begin
       hitMadPrint68 = 0;
    end
  end
end


string linebuf69 = "";
logic hitMadPrint69 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc69_inst_done && ((spc69_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint69 = 1;
       linebuf69 = {linebuf69, spc69_phy_pc_w[8:1]};
       if (spc69_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 69, linebuf69);
          linebuf69 = "";
       end
    end else begin
       hitMadPrint69 = 0;
    end
  end
end


string linebuf70 = "";
logic hitMadPrint70 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc70_inst_done && ((spc70_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint70 = 1;
       linebuf70 = {linebuf70, spc70_phy_pc_w[8:1]};
       if (spc70_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 70, linebuf70);
          linebuf70 = "";
       end
    end else begin
       hitMadPrint70 = 0;
    end
  end
end


string linebuf71 = "";
logic hitMadPrint71 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc71_inst_done && ((spc71_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint71 = 1;
       linebuf71 = {linebuf71, spc71_phy_pc_w[8:1]};
       if (spc71_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 71, linebuf71);
          linebuf71 = "";
       end
    end else begin
       hitMadPrint71 = 0;
    end
  end
end


string linebuf72 = "";
logic hitMadPrint72 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc72_inst_done && ((spc72_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint72 = 1;
       linebuf72 = {linebuf72, spc72_phy_pc_w[8:1]};
       if (spc72_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 72, linebuf72);
          linebuf72 = "";
       end
    end else begin
       hitMadPrint72 = 0;
    end
  end
end


string linebuf73 = "";
logic hitMadPrint73 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc73_inst_done && ((spc73_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint73 = 1;
       linebuf73 = {linebuf73, spc73_phy_pc_w[8:1]};
       if (spc73_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 73, linebuf73);
          linebuf73 = "";
       end
    end else begin
       hitMadPrint73 = 0;
    end
  end
end


string linebuf74 = "";
logic hitMadPrint74 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc74_inst_done && ((spc74_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint74 = 1;
       linebuf74 = {linebuf74, spc74_phy_pc_w[8:1]};
       if (spc74_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 74, linebuf74);
          linebuf74 = "";
       end
    end else begin
       hitMadPrint74 = 0;
    end
  end
end


string linebuf75 = "";
logic hitMadPrint75 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc75_inst_done && ((spc75_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint75 = 1;
       linebuf75 = {linebuf75, spc75_phy_pc_w[8:1]};
       if (spc75_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 75, linebuf75);
          linebuf75 = "";
       end
    end else begin
       hitMadPrint75 = 0;
    end
  end
end


string linebuf76 = "";
logic hitMadPrint76 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc76_inst_done && ((spc76_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint76 = 1;
       linebuf76 = {linebuf76, spc76_phy_pc_w[8:1]};
       if (spc76_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 76, linebuf76);
          linebuf76 = "";
       end
    end else begin
       hitMadPrint76 = 0;
    end
  end
end


string linebuf77 = "";
logic hitMadPrint77 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc77_inst_done && ((spc77_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint77 = 1;
       linebuf77 = {linebuf77, spc77_phy_pc_w[8:1]};
       if (spc77_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 77, linebuf77);
          linebuf77 = "";
       end
    end else begin
       hitMadPrint77 = 0;
    end
  end
end


string linebuf78 = "";
logic hitMadPrint78 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc78_inst_done && ((spc78_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint78 = 1;
       linebuf78 = {linebuf78, spc78_phy_pc_w[8:1]};
       if (spc78_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 78, linebuf78);
          linebuf78 = "";
       end
    end else begin
       hitMadPrint78 = 0;
    end
  end
end


string linebuf79 = "";
logic hitMadPrint79 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc79_inst_done && ((spc79_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint79 = 1;
       linebuf79 = {linebuf79, spc79_phy_pc_w[8:1]};
       if (spc79_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 79, linebuf79);
          linebuf79 = "";
       end
    end else begin
       hitMadPrint79 = 0;
    end
  end
end


string linebuf80 = "";
logic hitMadPrint80 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc80_inst_done && ((spc80_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint80 = 1;
       linebuf80 = {linebuf80, spc80_phy_pc_w[8:1]};
       if (spc80_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 80, linebuf80);
          linebuf80 = "";
       end
    end else begin
       hitMadPrint80 = 0;
    end
  end
end


string linebuf81 = "";
logic hitMadPrint81 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc81_inst_done && ((spc81_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint81 = 1;
       linebuf81 = {linebuf81, spc81_phy_pc_w[8:1]};
       if (spc81_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 81, linebuf81);
          linebuf81 = "";
       end
    end else begin
       hitMadPrint81 = 0;
    end
  end
end


string linebuf82 = "";
logic hitMadPrint82 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc82_inst_done && ((spc82_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint82 = 1;
       linebuf82 = {linebuf82, spc82_phy_pc_w[8:1]};
       if (spc82_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 82, linebuf82);
          linebuf82 = "";
       end
    end else begin
       hitMadPrint82 = 0;
    end
  end
end


string linebuf83 = "";
logic hitMadPrint83 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc83_inst_done && ((spc83_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint83 = 1;
       linebuf83 = {linebuf83, spc83_phy_pc_w[8:1]};
       if (spc83_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 83, linebuf83);
          linebuf83 = "";
       end
    end else begin
       hitMadPrint83 = 0;
    end
  end
end


string linebuf84 = "";
logic hitMadPrint84 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc84_inst_done && ((spc84_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint84 = 1;
       linebuf84 = {linebuf84, spc84_phy_pc_w[8:1]};
       if (spc84_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 84, linebuf84);
          linebuf84 = "";
       end
    end else begin
       hitMadPrint84 = 0;
    end
  end
end


string linebuf85 = "";
logic hitMadPrint85 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc85_inst_done && ((spc85_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint85 = 1;
       linebuf85 = {linebuf85, spc85_phy_pc_w[8:1]};
       if (spc85_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 85, linebuf85);
          linebuf85 = "";
       end
    end else begin
       hitMadPrint85 = 0;
    end
  end
end


string linebuf86 = "";
logic hitMadPrint86 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc86_inst_done && ((spc86_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint86 = 1;
       linebuf86 = {linebuf86, spc86_phy_pc_w[8:1]};
       if (spc86_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 86, linebuf86);
          linebuf86 = "";
       end
    end else begin
       hitMadPrint86 = 0;
    end
  end
end


string linebuf87 = "";
logic hitMadPrint87 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc87_inst_done && ((spc87_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint87 = 1;
       linebuf87 = {linebuf87, spc87_phy_pc_w[8:1]};
       if (spc87_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 87, linebuf87);
          linebuf87 = "";
       end
    end else begin
       hitMadPrint87 = 0;
    end
  end
end


string linebuf88 = "";
logic hitMadPrint88 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc88_inst_done && ((spc88_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint88 = 1;
       linebuf88 = {linebuf88, spc88_phy_pc_w[8:1]};
       if (spc88_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 88, linebuf88);
          linebuf88 = "";
       end
    end else begin
       hitMadPrint88 = 0;
    end
  end
end


string linebuf89 = "";
logic hitMadPrint89 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc89_inst_done && ((spc89_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint89 = 1;
       linebuf89 = {linebuf89, spc89_phy_pc_w[8:1]};
       if (spc89_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 89, linebuf89);
          linebuf89 = "";
       end
    end else begin
       hitMadPrint89 = 0;
    end
  end
end


string linebuf90 = "";
logic hitMadPrint90 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc90_inst_done && ((spc90_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint90 = 1;
       linebuf90 = {linebuf90, spc90_phy_pc_w[8:1]};
       if (spc90_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 90, linebuf90);
          linebuf90 = "";
       end
    end else begin
       hitMadPrint90 = 0;
    end
  end
end


string linebuf91 = "";
logic hitMadPrint91 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc91_inst_done && ((spc91_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint91 = 1;
       linebuf91 = {linebuf91, spc91_phy_pc_w[8:1]};
       if (spc91_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 91, linebuf91);
          linebuf91 = "";
       end
    end else begin
       hitMadPrint91 = 0;
    end
  end
end


string linebuf92 = "";
logic hitMadPrint92 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc92_inst_done && ((spc92_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint92 = 1;
       linebuf92 = {linebuf92, spc92_phy_pc_w[8:1]};
       if (spc92_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 92, linebuf92);
          linebuf92 = "";
       end
    end else begin
       hitMadPrint92 = 0;
    end
  end
end


string linebuf93 = "";
logic hitMadPrint93 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc93_inst_done && ((spc93_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint93 = 1;
       linebuf93 = {linebuf93, spc93_phy_pc_w[8:1]};
       if (spc93_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 93, linebuf93);
          linebuf93 = "";
       end
    end else begin
       hitMadPrint93 = 0;
    end
  end
end


string linebuf94 = "";
logic hitMadPrint94 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc94_inst_done && ((spc94_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint94 = 1;
       linebuf94 = {linebuf94, spc94_phy_pc_w[8:1]};
       if (spc94_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 94, linebuf94);
          linebuf94 = "";
       end
    end else begin
       hitMadPrint94 = 0;
    end
  end
end


string linebuf95 = "";
logic hitMadPrint95 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc95_inst_done && ((spc95_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint95 = 1;
       linebuf95 = {linebuf95, spc95_phy_pc_w[8:1]};
       if (spc95_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 95, linebuf95);
          linebuf95 = "";
       end
    end else begin
       hitMadPrint95 = 0;
    end
  end
end


string linebuf96 = "";
logic hitMadPrint96 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc96_inst_done && ((spc96_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint96 = 1;
       linebuf96 = {linebuf96, spc96_phy_pc_w[8:1]};
       if (spc96_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 96, linebuf96);
          linebuf96 = "";
       end
    end else begin
       hitMadPrint96 = 0;
    end
  end
end


string linebuf97 = "";
logic hitMadPrint97 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc97_inst_done && ((spc97_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint97 = 1;
       linebuf97 = {linebuf97, spc97_phy_pc_w[8:1]};
       if (spc97_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 97, linebuf97);
          linebuf97 = "";
       end
    end else begin
       hitMadPrint97 = 0;
    end
  end
end


string linebuf98 = "";
logic hitMadPrint98 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc98_inst_done && ((spc98_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint98 = 1;
       linebuf98 = {linebuf98, spc98_phy_pc_w[8:1]};
       if (spc98_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 98, linebuf98);
          linebuf98 = "";
       end
    end else begin
       hitMadPrint98 = 0;
    end
  end
end


string linebuf99 = "";
logic hitMadPrint99 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc99_inst_done && ((spc99_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint99 = 1;
       linebuf99 = {linebuf99, spc99_phy_pc_w[8:1]};
       if (spc99_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 99, linebuf99);
          linebuf99 = "";
       end
    end else begin
       hitMadPrint99 = 0;
    end
  end
end


string linebuf100 = "";
logic hitMadPrint100 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc100_inst_done && ((spc100_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint100 = 1;
       linebuf100 = {linebuf100, spc100_phy_pc_w[8:1]};
       if (spc100_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 100, linebuf100);
          linebuf100 = "";
       end
    end else begin
       hitMadPrint100 = 0;
    end
  end
end


string linebuf101 = "";
logic hitMadPrint101 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc101_inst_done && ((spc101_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint101 = 1;
       linebuf101 = {linebuf101, spc101_phy_pc_w[8:1]};
       if (spc101_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 101, linebuf101);
          linebuf101 = "";
       end
    end else begin
       hitMadPrint101 = 0;
    end
  end
end


string linebuf102 = "";
logic hitMadPrint102 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc102_inst_done && ((spc102_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint102 = 1;
       linebuf102 = {linebuf102, spc102_phy_pc_w[8:1]};
       if (spc102_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 102, linebuf102);
          linebuf102 = "";
       end
    end else begin
       hitMadPrint102 = 0;
    end
  end
end


string linebuf103 = "";
logic hitMadPrint103 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc103_inst_done && ((spc103_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint103 = 1;
       linebuf103 = {linebuf103, spc103_phy_pc_w[8:1]};
       if (spc103_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 103, linebuf103);
          linebuf103 = "";
       end
    end else begin
       hitMadPrint103 = 0;
    end
  end
end


string linebuf104 = "";
logic hitMadPrint104 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc104_inst_done && ((spc104_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint104 = 1;
       linebuf104 = {linebuf104, spc104_phy_pc_w[8:1]};
       if (spc104_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 104, linebuf104);
          linebuf104 = "";
       end
    end else begin
       hitMadPrint104 = 0;
    end
  end
end


string linebuf105 = "";
logic hitMadPrint105 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc105_inst_done && ((spc105_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint105 = 1;
       linebuf105 = {linebuf105, spc105_phy_pc_w[8:1]};
       if (spc105_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 105, linebuf105);
          linebuf105 = "";
       end
    end else begin
       hitMadPrint105 = 0;
    end
  end
end


string linebuf106 = "";
logic hitMadPrint106 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc106_inst_done && ((spc106_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint106 = 1;
       linebuf106 = {linebuf106, spc106_phy_pc_w[8:1]};
       if (spc106_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 106, linebuf106);
          linebuf106 = "";
       end
    end else begin
       hitMadPrint106 = 0;
    end
  end
end


string linebuf107 = "";
logic hitMadPrint107 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc107_inst_done && ((spc107_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint107 = 1;
       linebuf107 = {linebuf107, spc107_phy_pc_w[8:1]};
       if (spc107_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 107, linebuf107);
          linebuf107 = "";
       end
    end else begin
       hitMadPrint107 = 0;
    end
  end
end


string linebuf108 = "";
logic hitMadPrint108 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc108_inst_done && ((spc108_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint108 = 1;
       linebuf108 = {linebuf108, spc108_phy_pc_w[8:1]};
       if (spc108_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 108, linebuf108);
          linebuf108 = "";
       end
    end else begin
       hitMadPrint108 = 0;
    end
  end
end


string linebuf109 = "";
logic hitMadPrint109 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc109_inst_done && ((spc109_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint109 = 1;
       linebuf109 = {linebuf109, spc109_phy_pc_w[8:1]};
       if (spc109_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 109, linebuf109);
          linebuf109 = "";
       end
    end else begin
       hitMadPrint109 = 0;
    end
  end
end


string linebuf110 = "";
logic hitMadPrint110 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc110_inst_done && ((spc110_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint110 = 1;
       linebuf110 = {linebuf110, spc110_phy_pc_w[8:1]};
       if (spc110_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 110, linebuf110);
          linebuf110 = "";
       end
    end else begin
       hitMadPrint110 = 0;
    end
  end
end


string linebuf111 = "";
logic hitMadPrint111 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc111_inst_done && ((spc111_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint111 = 1;
       linebuf111 = {linebuf111, spc111_phy_pc_w[8:1]};
       if (spc111_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 111, linebuf111);
          linebuf111 = "";
       end
    end else begin
       hitMadPrint111 = 0;
    end
  end
end


string linebuf112 = "";
logic hitMadPrint112 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc112_inst_done && ((spc112_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint112 = 1;
       linebuf112 = {linebuf112, spc112_phy_pc_w[8:1]};
       if (spc112_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 112, linebuf112);
          linebuf112 = "";
       end
    end else begin
       hitMadPrint112 = 0;
    end
  end
end


string linebuf113 = "";
logic hitMadPrint113 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc113_inst_done && ((spc113_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint113 = 1;
       linebuf113 = {linebuf113, spc113_phy_pc_w[8:1]};
       if (spc113_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 113, linebuf113);
          linebuf113 = "";
       end
    end else begin
       hitMadPrint113 = 0;
    end
  end
end


string linebuf114 = "";
logic hitMadPrint114 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc114_inst_done && ((spc114_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint114 = 1;
       linebuf114 = {linebuf114, spc114_phy_pc_w[8:1]};
       if (spc114_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 114, linebuf114);
          linebuf114 = "";
       end
    end else begin
       hitMadPrint114 = 0;
    end
  end
end


string linebuf115 = "";
logic hitMadPrint115 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc115_inst_done && ((spc115_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint115 = 1;
       linebuf115 = {linebuf115, spc115_phy_pc_w[8:1]};
       if (spc115_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 115, linebuf115);
          linebuf115 = "";
       end
    end else begin
       hitMadPrint115 = 0;
    end
  end
end


string linebuf116 = "";
logic hitMadPrint116 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc116_inst_done && ((spc116_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint116 = 1;
       linebuf116 = {linebuf116, spc116_phy_pc_w[8:1]};
       if (spc116_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 116, linebuf116);
          linebuf116 = "";
       end
    end else begin
       hitMadPrint116 = 0;
    end
  end
end


string linebuf117 = "";
logic hitMadPrint117 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc117_inst_done && ((spc117_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint117 = 1;
       linebuf117 = {linebuf117, spc117_phy_pc_w[8:1]};
       if (spc117_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 117, linebuf117);
          linebuf117 = "";
       end
    end else begin
       hitMadPrint117 = 0;
    end
  end
end


string linebuf118 = "";
logic hitMadPrint118 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc118_inst_done && ((spc118_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint118 = 1;
       linebuf118 = {linebuf118, spc118_phy_pc_w[8:1]};
       if (spc118_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 118, linebuf118);
          linebuf118 = "";
       end
    end else begin
       hitMadPrint118 = 0;
    end
  end
end


string linebuf119 = "";
logic hitMadPrint119 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc119_inst_done && ((spc119_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint119 = 1;
       linebuf119 = {linebuf119, spc119_phy_pc_w[8:1]};
       if (spc119_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 119, linebuf119);
          linebuf119 = "";
       end
    end else begin
       hitMadPrint119 = 0;
    end
  end
end


string linebuf120 = "";
logic hitMadPrint120 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc120_inst_done && ((spc120_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint120 = 1;
       linebuf120 = {linebuf120, spc120_phy_pc_w[8:1]};
       if (spc120_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 120, linebuf120);
          linebuf120 = "";
       end
    end else begin
       hitMadPrint120 = 0;
    end
  end
end


string linebuf121 = "";
logic hitMadPrint121 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc121_inst_done && ((spc121_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint121 = 1;
       linebuf121 = {linebuf121, spc121_phy_pc_w[8:1]};
       if (spc121_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 121, linebuf121);
          linebuf121 = "";
       end
    end else begin
       hitMadPrint121 = 0;
    end
  end
end


string linebuf122 = "";
logic hitMadPrint122 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc122_inst_done && ((spc122_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint122 = 1;
       linebuf122 = {linebuf122, spc122_phy_pc_w[8:1]};
       if (spc122_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 122, linebuf122);
          linebuf122 = "";
       end
    end else begin
       hitMadPrint122 = 0;
    end
  end
end


string linebuf123 = "";
logic hitMadPrint123 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc123_inst_done && ((spc123_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint123 = 1;
       linebuf123 = {linebuf123, spc123_phy_pc_w[8:1]};
       if (spc123_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 123, linebuf123);
          linebuf123 = "";
       end
    end else begin
       hitMadPrint123 = 0;
    end
  end
end


string linebuf124 = "";
logic hitMadPrint124 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc124_inst_done && ((spc124_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint124 = 1;
       linebuf124 = {linebuf124, spc124_phy_pc_w[8:1]};
       if (spc124_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 124, linebuf124);
          linebuf124 = "";
       end
    end else begin
       hitMadPrint124 = 0;
    end
  end
end


string linebuf125 = "";
logic hitMadPrint125 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc125_inst_done && ((spc125_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint125 = 1;
       linebuf125 = {linebuf125, spc125_phy_pc_w[8:1]};
       if (spc125_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 125, linebuf125);
          linebuf125 = "";
       end
    end else begin
       hitMadPrint125 = 0;
    end
  end
end


string linebuf126 = "";
logic hitMadPrint126 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc126_inst_done && ((spc126_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint126 = 1;
       linebuf126 = {linebuf126, spc126_phy_pc_w[8:1]};
       if (spc126_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 126, linebuf126);
          linebuf126 = "";
       end
    end else begin
       hitMadPrint126 = 0;
    end
  end
end


string linebuf127 = "";
logic hitMadPrint127 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc127_inst_done && ((spc127_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint127 = 1;
       linebuf127 = {linebuf127, spc127_phy_pc_w[8:1]};
       if (spc127_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 127, linebuf127);
          linebuf127 = "";
       end
    end else begin
       hitMadPrint127 = 0;
    end
  end
end


string linebuf128 = "";
logic hitMadPrint128 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc128_inst_done && ((spc128_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint128 = 1;
       linebuf128 = {linebuf128, spc128_phy_pc_w[8:1]};
       if (spc128_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 128, linebuf128);
          linebuf128 = "";
       end
    end else begin
       hitMadPrint128 = 0;
    end
  end
end


string linebuf129 = "";
logic hitMadPrint129 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc129_inst_done && ((spc129_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint129 = 1;
       linebuf129 = {linebuf129, spc129_phy_pc_w[8:1]};
       if (spc129_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 129, linebuf129);
          linebuf129 = "";
       end
    end else begin
       hitMadPrint129 = 0;
    end
  end
end


string linebuf130 = "";
logic hitMadPrint130 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc130_inst_done && ((spc130_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint130 = 1;
       linebuf130 = {linebuf130, spc130_phy_pc_w[8:1]};
       if (spc130_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 130, linebuf130);
          linebuf130 = "";
       end
    end else begin
       hitMadPrint130 = 0;
    end
  end
end


string linebuf131 = "";
logic hitMadPrint131 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc131_inst_done && ((spc131_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint131 = 1;
       linebuf131 = {linebuf131, spc131_phy_pc_w[8:1]};
       if (spc131_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 131, linebuf131);
          linebuf131 = "";
       end
    end else begin
       hitMadPrint131 = 0;
    end
  end
end


string linebuf132 = "";
logic hitMadPrint132 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc132_inst_done && ((spc132_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint132 = 1;
       linebuf132 = {linebuf132, spc132_phy_pc_w[8:1]};
       if (spc132_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 132, linebuf132);
          linebuf132 = "";
       end
    end else begin
       hitMadPrint132 = 0;
    end
  end
end


string linebuf133 = "";
logic hitMadPrint133 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc133_inst_done && ((spc133_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint133 = 1;
       linebuf133 = {linebuf133, spc133_phy_pc_w[8:1]};
       if (spc133_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 133, linebuf133);
          linebuf133 = "";
       end
    end else begin
       hitMadPrint133 = 0;
    end
  end
end


string linebuf134 = "";
logic hitMadPrint134 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc134_inst_done && ((spc134_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint134 = 1;
       linebuf134 = {linebuf134, spc134_phy_pc_w[8:1]};
       if (spc134_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 134, linebuf134);
          linebuf134 = "";
       end
    end else begin
       hitMadPrint134 = 0;
    end
  end
end


string linebuf135 = "";
logic hitMadPrint135 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc135_inst_done && ((spc135_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint135 = 1;
       linebuf135 = {linebuf135, spc135_phy_pc_w[8:1]};
       if (spc135_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 135, linebuf135);
          linebuf135 = "";
       end
    end else begin
       hitMadPrint135 = 0;
    end
  end
end


string linebuf136 = "";
logic hitMadPrint136 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc136_inst_done && ((spc136_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint136 = 1;
       linebuf136 = {linebuf136, spc136_phy_pc_w[8:1]};
       if (spc136_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 136, linebuf136);
          linebuf136 = "";
       end
    end else begin
       hitMadPrint136 = 0;
    end
  end
end


string linebuf137 = "";
logic hitMadPrint137 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc137_inst_done && ((spc137_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint137 = 1;
       linebuf137 = {linebuf137, spc137_phy_pc_w[8:1]};
       if (spc137_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 137, linebuf137);
          linebuf137 = "";
       end
    end else begin
       hitMadPrint137 = 0;
    end
  end
end


string linebuf138 = "";
logic hitMadPrint138 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc138_inst_done && ((spc138_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint138 = 1;
       linebuf138 = {linebuf138, spc138_phy_pc_w[8:1]};
       if (spc138_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 138, linebuf138);
          linebuf138 = "";
       end
    end else begin
       hitMadPrint138 = 0;
    end
  end
end


string linebuf139 = "";
logic hitMadPrint139 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc139_inst_done && ((spc139_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint139 = 1;
       linebuf139 = {linebuf139, spc139_phy_pc_w[8:1]};
       if (spc139_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 139, linebuf139);
          linebuf139 = "";
       end
    end else begin
       hitMadPrint139 = 0;
    end
  end
end


string linebuf140 = "";
logic hitMadPrint140 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc140_inst_done && ((spc140_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint140 = 1;
       linebuf140 = {linebuf140, spc140_phy_pc_w[8:1]};
       if (spc140_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 140, linebuf140);
          linebuf140 = "";
       end
    end else begin
       hitMadPrint140 = 0;
    end
  end
end


string linebuf141 = "";
logic hitMadPrint141 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc141_inst_done && ((spc141_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint141 = 1;
       linebuf141 = {linebuf141, spc141_phy_pc_w[8:1]};
       if (spc141_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 141, linebuf141);
          linebuf141 = "";
       end
    end else begin
       hitMadPrint141 = 0;
    end
  end
end


string linebuf142 = "";
logic hitMadPrint142 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc142_inst_done && ((spc142_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint142 = 1;
       linebuf142 = {linebuf142, spc142_phy_pc_w[8:1]};
       if (spc142_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 142, linebuf142);
          linebuf142 = "";
       end
    end else begin
       hitMadPrint142 = 0;
    end
  end
end


string linebuf143 = "";
logic hitMadPrint143 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc143_inst_done && ((spc143_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint143 = 1;
       linebuf143 = {linebuf143, spc143_phy_pc_w[8:1]};
       if (spc143_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 143, linebuf143);
          linebuf143 = "";
       end
    end else begin
       hitMadPrint143 = 0;
    end
  end
end


string linebuf144 = "";
logic hitMadPrint144 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc144_inst_done && ((spc144_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint144 = 1;
       linebuf144 = {linebuf144, spc144_phy_pc_w[8:1]};
       if (spc144_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 144, linebuf144);
          linebuf144 = "";
       end
    end else begin
       hitMadPrint144 = 0;
    end
  end
end


string linebuf145 = "";
logic hitMadPrint145 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc145_inst_done && ((spc145_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint145 = 1;
       linebuf145 = {linebuf145, spc145_phy_pc_w[8:1]};
       if (spc145_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 145, linebuf145);
          linebuf145 = "";
       end
    end else begin
       hitMadPrint145 = 0;
    end
  end
end


string linebuf146 = "";
logic hitMadPrint146 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc146_inst_done && ((spc146_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint146 = 1;
       linebuf146 = {linebuf146, spc146_phy_pc_w[8:1]};
       if (spc146_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 146, linebuf146);
          linebuf146 = "";
       end
    end else begin
       hitMadPrint146 = 0;
    end
  end
end


string linebuf147 = "";
logic hitMadPrint147 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc147_inst_done && ((spc147_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint147 = 1;
       linebuf147 = {linebuf147, spc147_phy_pc_w[8:1]};
       if (spc147_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 147, linebuf147);
          linebuf147 = "";
       end
    end else begin
       hitMadPrint147 = 0;
    end
  end
end


string linebuf148 = "";
logic hitMadPrint148 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc148_inst_done && ((spc148_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint148 = 1;
       linebuf148 = {linebuf148, spc148_phy_pc_w[8:1]};
       if (spc148_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 148, linebuf148);
          linebuf148 = "";
       end
    end else begin
       hitMadPrint148 = 0;
    end
  end
end


string linebuf149 = "";
logic hitMadPrint149 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc149_inst_done && ((spc149_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint149 = 1;
       linebuf149 = {linebuf149, spc149_phy_pc_w[8:1]};
       if (spc149_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 149, linebuf149);
          linebuf149 = "";
       end
    end else begin
       hitMadPrint149 = 0;
    end
  end
end


string linebuf150 = "";
logic hitMadPrint150 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc150_inst_done && ((spc150_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint150 = 1;
       linebuf150 = {linebuf150, spc150_phy_pc_w[8:1]};
       if (spc150_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 150, linebuf150);
          linebuf150 = "";
       end
    end else begin
       hitMadPrint150 = 0;
    end
  end
end


string linebuf151 = "";
logic hitMadPrint151 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc151_inst_done && ((spc151_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint151 = 1;
       linebuf151 = {linebuf151, spc151_phy_pc_w[8:1]};
       if (spc151_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 151, linebuf151);
          linebuf151 = "";
       end
    end else begin
       hitMadPrint151 = 0;
    end
  end
end


string linebuf152 = "";
logic hitMadPrint152 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc152_inst_done && ((spc152_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint152 = 1;
       linebuf152 = {linebuf152, spc152_phy_pc_w[8:1]};
       if (spc152_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 152, linebuf152);
          linebuf152 = "";
       end
    end else begin
       hitMadPrint152 = 0;
    end
  end
end


string linebuf153 = "";
logic hitMadPrint153 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc153_inst_done && ((spc153_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint153 = 1;
       linebuf153 = {linebuf153, spc153_phy_pc_w[8:1]};
       if (spc153_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 153, linebuf153);
          linebuf153 = "";
       end
    end else begin
       hitMadPrint153 = 0;
    end
  end
end


string linebuf154 = "";
logic hitMadPrint154 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc154_inst_done && ((spc154_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint154 = 1;
       linebuf154 = {linebuf154, spc154_phy_pc_w[8:1]};
       if (spc154_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 154, linebuf154);
          linebuf154 = "";
       end
    end else begin
       hitMadPrint154 = 0;
    end
  end
end


string linebuf155 = "";
logic hitMadPrint155 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc155_inst_done && ((spc155_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint155 = 1;
       linebuf155 = {linebuf155, spc155_phy_pc_w[8:1]};
       if (spc155_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 155, linebuf155);
          linebuf155 = "";
       end
    end else begin
       hitMadPrint155 = 0;
    end
  end
end


string linebuf156 = "";
logic hitMadPrint156 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc156_inst_done && ((spc156_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint156 = 1;
       linebuf156 = {linebuf156, spc156_phy_pc_w[8:1]};
       if (spc156_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 156, linebuf156);
          linebuf156 = "";
       end
    end else begin
       hitMadPrint156 = 0;
    end
  end
end


string linebuf157 = "";
logic hitMadPrint157 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc157_inst_done && ((spc157_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint157 = 1;
       linebuf157 = {linebuf157, spc157_phy_pc_w[8:1]};
       if (spc157_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 157, linebuf157);
          linebuf157 = "";
       end
    end else begin
       hitMadPrint157 = 0;
    end
  end
end


string linebuf158 = "";
logic hitMadPrint158 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc158_inst_done && ((spc158_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint158 = 1;
       linebuf158 = {linebuf158, spc158_phy_pc_w[8:1]};
       if (spc158_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 158, linebuf158);
          linebuf158 = "";
       end
    end else begin
       hitMadPrint158 = 0;
    end
  end
end


string linebuf159 = "";
logic hitMadPrint159 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc159_inst_done && ((spc159_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint159 = 1;
       linebuf159 = {linebuf159, spc159_phy_pc_w[8:1]};
       if (spc159_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 159, linebuf159);
          linebuf159 = "";
       end
    end else begin
       hitMadPrint159 = 0;
    end
  end
end


string linebuf160 = "";
logic hitMadPrint160 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc160_inst_done && ((spc160_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint160 = 1;
       linebuf160 = {linebuf160, spc160_phy_pc_w[8:1]};
       if (spc160_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 160, linebuf160);
          linebuf160 = "";
       end
    end else begin
       hitMadPrint160 = 0;
    end
  end
end


string linebuf161 = "";
logic hitMadPrint161 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc161_inst_done && ((spc161_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint161 = 1;
       linebuf161 = {linebuf161, spc161_phy_pc_w[8:1]};
       if (spc161_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 161, linebuf161);
          linebuf161 = "";
       end
    end else begin
       hitMadPrint161 = 0;
    end
  end
end


string linebuf162 = "";
logic hitMadPrint162 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc162_inst_done && ((spc162_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint162 = 1;
       linebuf162 = {linebuf162, spc162_phy_pc_w[8:1]};
       if (spc162_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 162, linebuf162);
          linebuf162 = "";
       end
    end else begin
       hitMadPrint162 = 0;
    end
  end
end


string linebuf163 = "";
logic hitMadPrint163 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc163_inst_done && ((spc163_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint163 = 1;
       linebuf163 = {linebuf163, spc163_phy_pc_w[8:1]};
       if (spc163_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 163, linebuf163);
          linebuf163 = "";
       end
    end else begin
       hitMadPrint163 = 0;
    end
  end
end


string linebuf164 = "";
logic hitMadPrint164 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc164_inst_done && ((spc164_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint164 = 1;
       linebuf164 = {linebuf164, spc164_phy_pc_w[8:1]};
       if (spc164_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 164, linebuf164);
          linebuf164 = "";
       end
    end else begin
       hitMadPrint164 = 0;
    end
  end
end


string linebuf165 = "";
logic hitMadPrint165 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc165_inst_done && ((spc165_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint165 = 1;
       linebuf165 = {linebuf165, spc165_phy_pc_w[8:1]};
       if (spc165_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 165, linebuf165);
          linebuf165 = "";
       end
    end else begin
       hitMadPrint165 = 0;
    end
  end
end


string linebuf166 = "";
logic hitMadPrint166 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc166_inst_done && ((spc166_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint166 = 1;
       linebuf166 = {linebuf166, spc166_phy_pc_w[8:1]};
       if (spc166_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 166, linebuf166);
          linebuf166 = "";
       end
    end else begin
       hitMadPrint166 = 0;
    end
  end
end


string linebuf167 = "";
logic hitMadPrint167 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc167_inst_done && ((spc167_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint167 = 1;
       linebuf167 = {linebuf167, spc167_phy_pc_w[8:1]};
       if (spc167_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 167, linebuf167);
          linebuf167 = "";
       end
    end else begin
       hitMadPrint167 = 0;
    end
  end
end


string linebuf168 = "";
logic hitMadPrint168 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc168_inst_done && ((spc168_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint168 = 1;
       linebuf168 = {linebuf168, spc168_phy_pc_w[8:1]};
       if (spc168_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 168, linebuf168);
          linebuf168 = "";
       end
    end else begin
       hitMadPrint168 = 0;
    end
  end
end


string linebuf169 = "";
logic hitMadPrint169 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc169_inst_done && ((spc169_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint169 = 1;
       linebuf169 = {linebuf169, spc169_phy_pc_w[8:1]};
       if (spc169_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 169, linebuf169);
          linebuf169 = "";
       end
    end else begin
       hitMadPrint169 = 0;
    end
  end
end


string linebuf170 = "";
logic hitMadPrint170 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc170_inst_done && ((spc170_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint170 = 1;
       linebuf170 = {linebuf170, spc170_phy_pc_w[8:1]};
       if (spc170_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 170, linebuf170);
          linebuf170 = "";
       end
    end else begin
       hitMadPrint170 = 0;
    end
  end
end


string linebuf171 = "";
logic hitMadPrint171 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc171_inst_done && ((spc171_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint171 = 1;
       linebuf171 = {linebuf171, spc171_phy_pc_w[8:1]};
       if (spc171_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 171, linebuf171);
          linebuf171 = "";
       end
    end else begin
       hitMadPrint171 = 0;
    end
  end
end


string linebuf172 = "";
logic hitMadPrint172 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc172_inst_done && ((spc172_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint172 = 1;
       linebuf172 = {linebuf172, spc172_phy_pc_w[8:1]};
       if (spc172_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 172, linebuf172);
          linebuf172 = "";
       end
    end else begin
       hitMadPrint172 = 0;
    end
  end
end


string linebuf173 = "";
logic hitMadPrint173 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc173_inst_done && ((spc173_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint173 = 1;
       linebuf173 = {linebuf173, spc173_phy_pc_w[8:1]};
       if (spc173_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 173, linebuf173);
          linebuf173 = "";
       end
    end else begin
       hitMadPrint173 = 0;
    end
  end
end


string linebuf174 = "";
logic hitMadPrint174 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc174_inst_done && ((spc174_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint174 = 1;
       linebuf174 = {linebuf174, spc174_phy_pc_w[8:1]};
       if (spc174_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 174, linebuf174);
          linebuf174 = "";
       end
    end else begin
       hitMadPrint174 = 0;
    end
  end
end


string linebuf175 = "";
logic hitMadPrint175 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc175_inst_done && ((spc175_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint175 = 1;
       linebuf175 = {linebuf175, spc175_phy_pc_w[8:1]};
       if (spc175_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 175, linebuf175);
          linebuf175 = "";
       end
    end else begin
       hitMadPrint175 = 0;
    end
  end
end


string linebuf176 = "";
logic hitMadPrint176 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc176_inst_done && ((spc176_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint176 = 1;
       linebuf176 = {linebuf176, spc176_phy_pc_w[8:1]};
       if (spc176_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 176, linebuf176);
          linebuf176 = "";
       end
    end else begin
       hitMadPrint176 = 0;
    end
  end
end


string linebuf177 = "";
logic hitMadPrint177 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc177_inst_done && ((spc177_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint177 = 1;
       linebuf177 = {linebuf177, spc177_phy_pc_w[8:1]};
       if (spc177_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 177, linebuf177);
          linebuf177 = "";
       end
    end else begin
       hitMadPrint177 = 0;
    end
  end
end


string linebuf178 = "";
logic hitMadPrint178 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc178_inst_done && ((spc178_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint178 = 1;
       linebuf178 = {linebuf178, spc178_phy_pc_w[8:1]};
       if (spc178_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 178, linebuf178);
          linebuf178 = "";
       end
    end else begin
       hitMadPrint178 = 0;
    end
  end
end


string linebuf179 = "";
logic hitMadPrint179 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc179_inst_done && ((spc179_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint179 = 1;
       linebuf179 = {linebuf179, spc179_phy_pc_w[8:1]};
       if (spc179_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 179, linebuf179);
          linebuf179 = "";
       end
    end else begin
       hitMadPrint179 = 0;
    end
  end
end


string linebuf180 = "";
logic hitMadPrint180 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc180_inst_done && ((spc180_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint180 = 1;
       linebuf180 = {linebuf180, spc180_phy_pc_w[8:1]};
       if (spc180_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 180, linebuf180);
          linebuf180 = "";
       end
    end else begin
       hitMadPrint180 = 0;
    end
  end
end


string linebuf181 = "";
logic hitMadPrint181 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc181_inst_done && ((spc181_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint181 = 1;
       linebuf181 = {linebuf181, spc181_phy_pc_w[8:1]};
       if (spc181_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 181, linebuf181);
          linebuf181 = "";
       end
    end else begin
       hitMadPrint181 = 0;
    end
  end
end


string linebuf182 = "";
logic hitMadPrint182 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc182_inst_done && ((spc182_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint182 = 1;
       linebuf182 = {linebuf182, spc182_phy_pc_w[8:1]};
       if (spc182_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 182, linebuf182);
          linebuf182 = "";
       end
    end else begin
       hitMadPrint182 = 0;
    end
  end
end


string linebuf183 = "";
logic hitMadPrint183 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc183_inst_done && ((spc183_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint183 = 1;
       linebuf183 = {linebuf183, spc183_phy_pc_w[8:1]};
       if (spc183_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 183, linebuf183);
          linebuf183 = "";
       end
    end else begin
       hitMadPrint183 = 0;
    end
  end
end


string linebuf184 = "";
logic hitMadPrint184 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc184_inst_done && ((spc184_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint184 = 1;
       linebuf184 = {linebuf184, spc184_phy_pc_w[8:1]};
       if (spc184_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 184, linebuf184);
          linebuf184 = "";
       end
    end else begin
       hitMadPrint184 = 0;
    end
  end
end


string linebuf185 = "";
logic hitMadPrint185 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc185_inst_done && ((spc185_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint185 = 1;
       linebuf185 = {linebuf185, spc185_phy_pc_w[8:1]};
       if (spc185_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 185, linebuf185);
          linebuf185 = "";
       end
    end else begin
       hitMadPrint185 = 0;
    end
  end
end


string linebuf186 = "";
logic hitMadPrint186 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc186_inst_done && ((spc186_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint186 = 1;
       linebuf186 = {linebuf186, spc186_phy_pc_w[8:1]};
       if (spc186_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 186, linebuf186);
          linebuf186 = "";
       end
    end else begin
       hitMadPrint186 = 0;
    end
  end
end


string linebuf187 = "";
logic hitMadPrint187 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc187_inst_done && ((spc187_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint187 = 1;
       linebuf187 = {linebuf187, spc187_phy_pc_w[8:1]};
       if (spc187_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 187, linebuf187);
          linebuf187 = "";
       end
    end else begin
       hitMadPrint187 = 0;
    end
  end
end


string linebuf188 = "";
logic hitMadPrint188 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc188_inst_done && ((spc188_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint188 = 1;
       linebuf188 = {linebuf188, spc188_phy_pc_w[8:1]};
       if (spc188_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 188, linebuf188);
          linebuf188 = "";
       end
    end else begin
       hitMadPrint188 = 0;
    end
  end
end


string linebuf189 = "";
logic hitMadPrint189 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc189_inst_done && ((spc189_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint189 = 1;
       linebuf189 = {linebuf189, spc189_phy_pc_w[8:1]};
       if (spc189_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 189, linebuf189);
          linebuf189 = "";
       end
    end else begin
       hitMadPrint189 = 0;
    end
  end
end


string linebuf190 = "";
logic hitMadPrint190 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc190_inst_done && ((spc190_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint190 = 1;
       linebuf190 = {linebuf190, spc190_phy_pc_w[8:1]};
       if (spc190_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 190, linebuf190);
          linebuf190 = "";
       end
    end else begin
       hitMadPrint190 = 0;
    end
  end
end


string linebuf191 = "";
logic hitMadPrint191 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc191_inst_done && ((spc191_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint191 = 1;
       linebuf191 = {linebuf191, spc191_phy_pc_w[8:1]};
       if (spc191_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 191, linebuf191);
          linebuf191 = "";
       end
    end else begin
       hitMadPrint191 = 0;
    end
  end
end


string linebuf192 = "";
logic hitMadPrint192 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc192_inst_done && ((spc192_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint192 = 1;
       linebuf192 = {linebuf192, spc192_phy_pc_w[8:1]};
       if (spc192_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 192, linebuf192);
          linebuf192 = "";
       end
    end else begin
       hitMadPrint192 = 0;
    end
  end
end


string linebuf193 = "";
logic hitMadPrint193 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc193_inst_done && ((spc193_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint193 = 1;
       linebuf193 = {linebuf193, spc193_phy_pc_w[8:1]};
       if (spc193_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 193, linebuf193);
          linebuf193 = "";
       end
    end else begin
       hitMadPrint193 = 0;
    end
  end
end


string linebuf194 = "";
logic hitMadPrint194 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc194_inst_done && ((spc194_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint194 = 1;
       linebuf194 = {linebuf194, spc194_phy_pc_w[8:1]};
       if (spc194_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 194, linebuf194);
          linebuf194 = "";
       end
    end else begin
       hitMadPrint194 = 0;
    end
  end
end


string linebuf195 = "";
logic hitMadPrint195 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc195_inst_done && ((spc195_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint195 = 1;
       linebuf195 = {linebuf195, spc195_phy_pc_w[8:1]};
       if (spc195_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 195, linebuf195);
          linebuf195 = "";
       end
    end else begin
       hitMadPrint195 = 0;
    end
  end
end


string linebuf196 = "";
logic hitMadPrint196 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc196_inst_done && ((spc196_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint196 = 1;
       linebuf196 = {linebuf196, spc196_phy_pc_w[8:1]};
       if (spc196_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 196, linebuf196);
          linebuf196 = "";
       end
    end else begin
       hitMadPrint196 = 0;
    end
  end
end


string linebuf197 = "";
logic hitMadPrint197 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc197_inst_done && ((spc197_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint197 = 1;
       linebuf197 = {linebuf197, spc197_phy_pc_w[8:1]};
       if (spc197_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 197, linebuf197);
          linebuf197 = "";
       end
    end else begin
       hitMadPrint197 = 0;
    end
  end
end


string linebuf198 = "";
logic hitMadPrint198 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc198_inst_done && ((spc198_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint198 = 1;
       linebuf198 = {linebuf198, spc198_phy_pc_w[8:1]};
       if (spc198_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 198, linebuf198);
          linebuf198 = "";
       end
    end else begin
       hitMadPrint198 = 0;
    end
  end
end


string linebuf199 = "";
logic hitMadPrint199 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc199_inst_done && ((spc199_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint199 = 1;
       linebuf199 = {linebuf199, spc199_phy_pc_w[8:1]};
       if (spc199_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 199, linebuf199);
          linebuf199 = "";
       end
    end else begin
       hitMadPrint199 = 0;
    end
  end
end


string linebuf200 = "";
logic hitMadPrint200 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc200_inst_done && ((spc200_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint200 = 1;
       linebuf200 = {linebuf200, spc200_phy_pc_w[8:1]};
       if (spc200_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 200, linebuf200);
          linebuf200 = "";
       end
    end else begin
       hitMadPrint200 = 0;
    end
  end
end


string linebuf201 = "";
logic hitMadPrint201 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc201_inst_done && ((spc201_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint201 = 1;
       linebuf201 = {linebuf201, spc201_phy_pc_w[8:1]};
       if (spc201_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 201, linebuf201);
          linebuf201 = "";
       end
    end else begin
       hitMadPrint201 = 0;
    end
  end
end


string linebuf202 = "";
logic hitMadPrint202 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc202_inst_done && ((spc202_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint202 = 1;
       linebuf202 = {linebuf202, spc202_phy_pc_w[8:1]};
       if (spc202_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 202, linebuf202);
          linebuf202 = "";
       end
    end else begin
       hitMadPrint202 = 0;
    end
  end
end


string linebuf203 = "";
logic hitMadPrint203 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc203_inst_done && ((spc203_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint203 = 1;
       linebuf203 = {linebuf203, spc203_phy_pc_w[8:1]};
       if (spc203_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 203, linebuf203);
          linebuf203 = "";
       end
    end else begin
       hitMadPrint203 = 0;
    end
  end
end


string linebuf204 = "";
logic hitMadPrint204 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc204_inst_done && ((spc204_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint204 = 1;
       linebuf204 = {linebuf204, spc204_phy_pc_w[8:1]};
       if (spc204_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 204, linebuf204);
          linebuf204 = "";
       end
    end else begin
       hitMadPrint204 = 0;
    end
  end
end


string linebuf205 = "";
logic hitMadPrint205 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc205_inst_done && ((spc205_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint205 = 1;
       linebuf205 = {linebuf205, spc205_phy_pc_w[8:1]};
       if (spc205_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 205, linebuf205);
          linebuf205 = "";
       end
    end else begin
       hitMadPrint205 = 0;
    end
  end
end


string linebuf206 = "";
logic hitMadPrint206 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc206_inst_done && ((spc206_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint206 = 1;
       linebuf206 = {linebuf206, spc206_phy_pc_w[8:1]};
       if (spc206_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 206, linebuf206);
          linebuf206 = "";
       end
    end else begin
       hitMadPrint206 = 0;
    end
  end
end


string linebuf207 = "";
logic hitMadPrint207 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc207_inst_done && ((spc207_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint207 = 1;
       linebuf207 = {linebuf207, spc207_phy_pc_w[8:1]};
       if (spc207_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 207, linebuf207);
          linebuf207 = "";
       end
    end else begin
       hitMadPrint207 = 0;
    end
  end
end


string linebuf208 = "";
logic hitMadPrint208 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc208_inst_done && ((spc208_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint208 = 1;
       linebuf208 = {linebuf208, spc208_phy_pc_w[8:1]};
       if (spc208_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 208, linebuf208);
          linebuf208 = "";
       end
    end else begin
       hitMadPrint208 = 0;
    end
  end
end


string linebuf209 = "";
logic hitMadPrint209 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc209_inst_done && ((spc209_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint209 = 1;
       linebuf209 = {linebuf209, spc209_phy_pc_w[8:1]};
       if (spc209_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 209, linebuf209);
          linebuf209 = "";
       end
    end else begin
       hitMadPrint209 = 0;
    end
  end
end


string linebuf210 = "";
logic hitMadPrint210 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc210_inst_done && ((spc210_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint210 = 1;
       linebuf210 = {linebuf210, spc210_phy_pc_w[8:1]};
       if (spc210_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 210, linebuf210);
          linebuf210 = "";
       end
    end else begin
       hitMadPrint210 = 0;
    end
  end
end


string linebuf211 = "";
logic hitMadPrint211 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc211_inst_done && ((spc211_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint211 = 1;
       linebuf211 = {linebuf211, spc211_phy_pc_w[8:1]};
       if (spc211_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 211, linebuf211);
          linebuf211 = "";
       end
    end else begin
       hitMadPrint211 = 0;
    end
  end
end


string linebuf212 = "";
logic hitMadPrint212 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc212_inst_done && ((spc212_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint212 = 1;
       linebuf212 = {linebuf212, spc212_phy_pc_w[8:1]};
       if (spc212_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 212, linebuf212);
          linebuf212 = "";
       end
    end else begin
       hitMadPrint212 = 0;
    end
  end
end


string linebuf213 = "";
logic hitMadPrint213 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc213_inst_done && ((spc213_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint213 = 1;
       linebuf213 = {linebuf213, spc213_phy_pc_w[8:1]};
       if (spc213_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 213, linebuf213);
          linebuf213 = "";
       end
    end else begin
       hitMadPrint213 = 0;
    end
  end
end


string linebuf214 = "";
logic hitMadPrint214 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc214_inst_done && ((spc214_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint214 = 1;
       linebuf214 = {linebuf214, spc214_phy_pc_w[8:1]};
       if (spc214_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 214, linebuf214);
          linebuf214 = "";
       end
    end else begin
       hitMadPrint214 = 0;
    end
  end
end


string linebuf215 = "";
logic hitMadPrint215 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc215_inst_done && ((spc215_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint215 = 1;
       linebuf215 = {linebuf215, spc215_phy_pc_w[8:1]};
       if (spc215_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 215, linebuf215);
          linebuf215 = "";
       end
    end else begin
       hitMadPrint215 = 0;
    end
  end
end


string linebuf216 = "";
logic hitMadPrint216 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc216_inst_done && ((spc216_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint216 = 1;
       linebuf216 = {linebuf216, spc216_phy_pc_w[8:1]};
       if (spc216_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 216, linebuf216);
          linebuf216 = "";
       end
    end else begin
       hitMadPrint216 = 0;
    end
  end
end


string linebuf217 = "";
logic hitMadPrint217 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc217_inst_done && ((spc217_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint217 = 1;
       linebuf217 = {linebuf217, spc217_phy_pc_w[8:1]};
       if (spc217_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 217, linebuf217);
          linebuf217 = "";
       end
    end else begin
       hitMadPrint217 = 0;
    end
  end
end


string linebuf218 = "";
logic hitMadPrint218 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc218_inst_done && ((spc218_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint218 = 1;
       linebuf218 = {linebuf218, spc218_phy_pc_w[8:1]};
       if (spc218_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 218, linebuf218);
          linebuf218 = "";
       end
    end else begin
       hitMadPrint218 = 0;
    end
  end
end


string linebuf219 = "";
logic hitMadPrint219 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc219_inst_done && ((spc219_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint219 = 1;
       linebuf219 = {linebuf219, spc219_phy_pc_w[8:1]};
       if (spc219_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 219, linebuf219);
          linebuf219 = "";
       end
    end else begin
       hitMadPrint219 = 0;
    end
  end
end


string linebuf220 = "";
logic hitMadPrint220 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc220_inst_done && ((spc220_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint220 = 1;
       linebuf220 = {linebuf220, spc220_phy_pc_w[8:1]};
       if (spc220_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 220, linebuf220);
          linebuf220 = "";
       end
    end else begin
       hitMadPrint220 = 0;
    end
  end
end


string linebuf221 = "";
logic hitMadPrint221 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc221_inst_done && ((spc221_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint221 = 1;
       linebuf221 = {linebuf221, spc221_phy_pc_w[8:1]};
       if (spc221_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 221, linebuf221);
          linebuf221 = "";
       end
    end else begin
       hitMadPrint221 = 0;
    end
  end
end


string linebuf222 = "";
logic hitMadPrint222 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc222_inst_done && ((spc222_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint222 = 1;
       linebuf222 = {linebuf222, spc222_phy_pc_w[8:1]};
       if (spc222_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 222, linebuf222);
          linebuf222 = "";
       end
    end else begin
       hitMadPrint222 = 0;
    end
  end
end


string linebuf223 = "";
logic hitMadPrint223 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc223_inst_done && ((spc223_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint223 = 1;
       linebuf223 = {linebuf223, spc223_phy_pc_w[8:1]};
       if (spc223_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 223, linebuf223);
          linebuf223 = "";
       end
    end else begin
       hitMadPrint223 = 0;
    end
  end
end


string linebuf224 = "";
logic hitMadPrint224 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc224_inst_done && ((spc224_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint224 = 1;
       linebuf224 = {linebuf224, spc224_phy_pc_w[8:1]};
       if (spc224_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 224, linebuf224);
          linebuf224 = "";
       end
    end else begin
       hitMadPrint224 = 0;
    end
  end
end


string linebuf225 = "";
logic hitMadPrint225 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc225_inst_done && ((spc225_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint225 = 1;
       linebuf225 = {linebuf225, spc225_phy_pc_w[8:1]};
       if (spc225_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 225, linebuf225);
          linebuf225 = "";
       end
    end else begin
       hitMadPrint225 = 0;
    end
  end
end


string linebuf226 = "";
logic hitMadPrint226 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc226_inst_done && ((spc226_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint226 = 1;
       linebuf226 = {linebuf226, spc226_phy_pc_w[8:1]};
       if (spc226_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 226, linebuf226);
          linebuf226 = "";
       end
    end else begin
       hitMadPrint226 = 0;
    end
  end
end


string linebuf227 = "";
logic hitMadPrint227 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc227_inst_done && ((spc227_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint227 = 1;
       linebuf227 = {linebuf227, spc227_phy_pc_w[8:1]};
       if (spc227_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 227, linebuf227);
          linebuf227 = "";
       end
    end else begin
       hitMadPrint227 = 0;
    end
  end
end


string linebuf228 = "";
logic hitMadPrint228 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc228_inst_done && ((spc228_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint228 = 1;
       linebuf228 = {linebuf228, spc228_phy_pc_w[8:1]};
       if (spc228_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 228, linebuf228);
          linebuf228 = "";
       end
    end else begin
       hitMadPrint228 = 0;
    end
  end
end


string linebuf229 = "";
logic hitMadPrint229 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc229_inst_done && ((spc229_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint229 = 1;
       linebuf229 = {linebuf229, spc229_phy_pc_w[8:1]};
       if (spc229_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 229, linebuf229);
          linebuf229 = "";
       end
    end else begin
       hitMadPrint229 = 0;
    end
  end
end


string linebuf230 = "";
logic hitMadPrint230 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc230_inst_done && ((spc230_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint230 = 1;
       linebuf230 = {linebuf230, spc230_phy_pc_w[8:1]};
       if (spc230_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 230, linebuf230);
          linebuf230 = "";
       end
    end else begin
       hitMadPrint230 = 0;
    end
  end
end


string linebuf231 = "";
logic hitMadPrint231 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc231_inst_done && ((spc231_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint231 = 1;
       linebuf231 = {linebuf231, spc231_phy_pc_w[8:1]};
       if (spc231_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 231, linebuf231);
          linebuf231 = "";
       end
    end else begin
       hitMadPrint231 = 0;
    end
  end
end


string linebuf232 = "";
logic hitMadPrint232 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc232_inst_done && ((spc232_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint232 = 1;
       linebuf232 = {linebuf232, spc232_phy_pc_w[8:1]};
       if (spc232_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 232, linebuf232);
          linebuf232 = "";
       end
    end else begin
       hitMadPrint232 = 0;
    end
  end
end


string linebuf233 = "";
logic hitMadPrint233 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc233_inst_done && ((spc233_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint233 = 1;
       linebuf233 = {linebuf233, spc233_phy_pc_w[8:1]};
       if (spc233_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 233, linebuf233);
          linebuf233 = "";
       end
    end else begin
       hitMadPrint233 = 0;
    end
  end
end


string linebuf234 = "";
logic hitMadPrint234 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc234_inst_done && ((spc234_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint234 = 1;
       linebuf234 = {linebuf234, spc234_phy_pc_w[8:1]};
       if (spc234_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 234, linebuf234);
          linebuf234 = "";
       end
    end else begin
       hitMadPrint234 = 0;
    end
  end
end


string linebuf235 = "";
logic hitMadPrint235 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc235_inst_done && ((spc235_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint235 = 1;
       linebuf235 = {linebuf235, spc235_phy_pc_w[8:1]};
       if (spc235_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 235, linebuf235);
          linebuf235 = "";
       end
    end else begin
       hitMadPrint235 = 0;
    end
  end
end


string linebuf236 = "";
logic hitMadPrint236 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc236_inst_done && ((spc236_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint236 = 1;
       linebuf236 = {linebuf236, spc236_phy_pc_w[8:1]};
       if (spc236_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 236, linebuf236);
          linebuf236 = "";
       end
    end else begin
       hitMadPrint236 = 0;
    end
  end
end


string linebuf237 = "";
logic hitMadPrint237 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc237_inst_done && ((spc237_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint237 = 1;
       linebuf237 = {linebuf237, spc237_phy_pc_w[8:1]};
       if (spc237_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 237, linebuf237);
          linebuf237 = "";
       end
    end else begin
       hitMadPrint237 = 0;
    end
  end
end


string linebuf238 = "";
logic hitMadPrint238 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc238_inst_done && ((spc238_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint238 = 1;
       linebuf238 = {linebuf238, spc238_phy_pc_w[8:1]};
       if (spc238_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 238, linebuf238);
          linebuf238 = "";
       end
    end else begin
       hitMadPrint238 = 0;
    end
  end
end


string linebuf239 = "";
logic hitMadPrint239 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc239_inst_done && ((spc239_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint239 = 1;
       linebuf239 = {linebuf239, spc239_phy_pc_w[8:1]};
       if (spc239_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 239, linebuf239);
          linebuf239 = "";
       end
    end else begin
       hitMadPrint239 = 0;
    end
  end
end


string linebuf240 = "";
logic hitMadPrint240 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc240_inst_done && ((spc240_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint240 = 1;
       linebuf240 = {linebuf240, spc240_phy_pc_w[8:1]};
       if (spc240_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 240, linebuf240);
          linebuf240 = "";
       end
    end else begin
       hitMadPrint240 = 0;
    end
  end
end


string linebuf241 = "";
logic hitMadPrint241 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc241_inst_done && ((spc241_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint241 = 1;
       linebuf241 = {linebuf241, spc241_phy_pc_w[8:1]};
       if (spc241_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 241, linebuf241);
          linebuf241 = "";
       end
    end else begin
       hitMadPrint241 = 0;
    end
  end
end


string linebuf242 = "";
logic hitMadPrint242 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc242_inst_done && ((spc242_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint242 = 1;
       linebuf242 = {linebuf242, spc242_phy_pc_w[8:1]};
       if (spc242_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 242, linebuf242);
          linebuf242 = "";
       end
    end else begin
       hitMadPrint242 = 0;
    end
  end
end


string linebuf243 = "";
logic hitMadPrint243 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc243_inst_done && ((spc243_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint243 = 1;
       linebuf243 = {linebuf243, spc243_phy_pc_w[8:1]};
       if (spc243_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 243, linebuf243);
          linebuf243 = "";
       end
    end else begin
       hitMadPrint243 = 0;
    end
  end
end


string linebuf244 = "";
logic hitMadPrint244 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc244_inst_done && ((spc244_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint244 = 1;
       linebuf244 = {linebuf244, spc244_phy_pc_w[8:1]};
       if (spc244_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 244, linebuf244);
          linebuf244 = "";
       end
    end else begin
       hitMadPrint244 = 0;
    end
  end
end


string linebuf245 = "";
logic hitMadPrint245 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc245_inst_done && ((spc245_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint245 = 1;
       linebuf245 = {linebuf245, spc245_phy_pc_w[8:1]};
       if (spc245_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 245, linebuf245);
          linebuf245 = "";
       end
    end else begin
       hitMadPrint245 = 0;
    end
  end
end


string linebuf246 = "";
logic hitMadPrint246 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc246_inst_done && ((spc246_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint246 = 1;
       linebuf246 = {linebuf246, spc246_phy_pc_w[8:1]};
       if (spc246_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 246, linebuf246);
          linebuf246 = "";
       end
    end else begin
       hitMadPrint246 = 0;
    end
  end
end


string linebuf247 = "";
logic hitMadPrint247 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc247_inst_done && ((spc247_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint247 = 1;
       linebuf247 = {linebuf247, spc247_phy_pc_w[8:1]};
       if (spc247_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 247, linebuf247);
          linebuf247 = "";
       end
    end else begin
       hitMadPrint247 = 0;
    end
  end
end


string linebuf248 = "";
logic hitMadPrint248 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc248_inst_done && ((spc248_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint248 = 1;
       linebuf248 = {linebuf248, spc248_phy_pc_w[8:1]};
       if (spc248_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 248, linebuf248);
          linebuf248 = "";
       end
    end else begin
       hitMadPrint248 = 0;
    end
  end
end


string linebuf249 = "";
logic hitMadPrint249 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc249_inst_done && ((spc249_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint249 = 1;
       linebuf249 = {linebuf249, spc249_phy_pc_w[8:1]};
       if (spc249_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 249, linebuf249);
          linebuf249 = "";
       end
    end else begin
       hitMadPrint249 = 0;
    end
  end
end


string linebuf250 = "";
logic hitMadPrint250 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc250_inst_done && ((spc250_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint250 = 1;
       linebuf250 = {linebuf250, spc250_phy_pc_w[8:1]};
       if (spc250_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 250, linebuf250);
          linebuf250 = "";
       end
    end else begin
       hitMadPrint250 = 0;
    end
  end
end


string linebuf251 = "";
logic hitMadPrint251 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc251_inst_done && ((spc251_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint251 = 1;
       linebuf251 = {linebuf251, spc251_phy_pc_w[8:1]};
       if (spc251_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 251, linebuf251);
          linebuf251 = "";
       end
    end else begin
       hitMadPrint251 = 0;
    end
  end
end


string linebuf252 = "";
logic hitMadPrint252 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc252_inst_done && ((spc252_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint252 = 1;
       linebuf252 = {linebuf252, spc252_phy_pc_w[8:1]};
       if (spc252_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 252, linebuf252);
          linebuf252 = "";
       end
    end else begin
       hitMadPrint252 = 0;
    end
  end
end


string linebuf253 = "";
logic hitMadPrint253 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc253_inst_done && ((spc253_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint253 = 1;
       linebuf253 = {linebuf253, spc253_phy_pc_w[8:1]};
       if (spc253_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 253, linebuf253);
          linebuf253 = "";
       end
    end else begin
       hitMadPrint253 = 0;
    end
  end
end


string linebuf254 = "";
logic hitMadPrint254 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc254_inst_done && ((spc254_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint254 = 1;
       linebuf254 = {linebuf254, spc254_phy_pc_w[8:1]};
       if (spc254_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 254, linebuf254);
          linebuf254 = "";
       end
    end else begin
       hitMadPrint254 = 0;
    end
  end
end


string linebuf255 = "";
logic hitMadPrint255 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc255_inst_done && ((spc255_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint255 = 1;
       linebuf255 = {linebuf255, spc255_phy_pc_w[8:1]};
       if (spc255_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 255, linebuf255);
          linebuf255 = "";
       end
    end else begin
       hitMadPrint255 = 0;
    end
  end
end


string linebuf256 = "";
logic hitMadPrint256 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc256_inst_done && ((spc256_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint256 = 1;
       linebuf256 = {linebuf256, spc256_phy_pc_w[8:1]};
       if (spc256_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 256, linebuf256);
          linebuf256 = "";
       end
    end else begin
       hitMadPrint256 = 0;
    end
  end
end


string linebuf257 = "";
logic hitMadPrint257 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc257_inst_done && ((spc257_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint257 = 1;
       linebuf257 = {linebuf257, spc257_phy_pc_w[8:1]};
       if (spc257_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 257, linebuf257);
          linebuf257 = "";
       end
    end else begin
       hitMadPrint257 = 0;
    end
  end
end


string linebuf258 = "";
logic hitMadPrint258 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc258_inst_done && ((spc258_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint258 = 1;
       linebuf258 = {linebuf258, spc258_phy_pc_w[8:1]};
       if (spc258_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 258, linebuf258);
          linebuf258 = "";
       end
    end else begin
       hitMadPrint258 = 0;
    end
  end
end


string linebuf259 = "";
logic hitMadPrint259 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc259_inst_done && ((spc259_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint259 = 1;
       linebuf259 = {linebuf259, spc259_phy_pc_w[8:1]};
       if (spc259_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 259, linebuf259);
          linebuf259 = "";
       end
    end else begin
       hitMadPrint259 = 0;
    end
  end
end


string linebuf260 = "";
logic hitMadPrint260 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc260_inst_done && ((spc260_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint260 = 1;
       linebuf260 = {linebuf260, spc260_phy_pc_w[8:1]};
       if (spc260_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 260, linebuf260);
          linebuf260 = "";
       end
    end else begin
       hitMadPrint260 = 0;
    end
  end
end


string linebuf261 = "";
logic hitMadPrint261 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc261_inst_done && ((spc261_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint261 = 1;
       linebuf261 = {linebuf261, spc261_phy_pc_w[8:1]};
       if (spc261_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 261, linebuf261);
          linebuf261 = "";
       end
    end else begin
       hitMadPrint261 = 0;
    end
  end
end


string linebuf262 = "";
logic hitMadPrint262 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc262_inst_done && ((spc262_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint262 = 1;
       linebuf262 = {linebuf262, spc262_phy_pc_w[8:1]};
       if (spc262_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 262, linebuf262);
          linebuf262 = "";
       end
    end else begin
       hitMadPrint262 = 0;
    end
  end
end


string linebuf263 = "";
logic hitMadPrint263 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc263_inst_done && ((spc263_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint263 = 1;
       linebuf263 = {linebuf263, spc263_phy_pc_w[8:1]};
       if (spc263_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 263, linebuf263);
          linebuf263 = "";
       end
    end else begin
       hitMadPrint263 = 0;
    end
  end
end


string linebuf264 = "";
logic hitMadPrint264 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc264_inst_done && ((spc264_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint264 = 1;
       linebuf264 = {linebuf264, spc264_phy_pc_w[8:1]};
       if (spc264_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 264, linebuf264);
          linebuf264 = "";
       end
    end else begin
       hitMadPrint264 = 0;
    end
  end
end


string linebuf265 = "";
logic hitMadPrint265 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc265_inst_done && ((spc265_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint265 = 1;
       linebuf265 = {linebuf265, spc265_phy_pc_w[8:1]};
       if (spc265_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 265, linebuf265);
          linebuf265 = "";
       end
    end else begin
       hitMadPrint265 = 0;
    end
  end
end


string linebuf266 = "";
logic hitMadPrint266 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc266_inst_done && ((spc266_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint266 = 1;
       linebuf266 = {linebuf266, spc266_phy_pc_w[8:1]};
       if (spc266_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 266, linebuf266);
          linebuf266 = "";
       end
    end else begin
       hitMadPrint266 = 0;
    end
  end
end


string linebuf267 = "";
logic hitMadPrint267 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc267_inst_done && ((spc267_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint267 = 1;
       linebuf267 = {linebuf267, spc267_phy_pc_w[8:1]};
       if (spc267_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 267, linebuf267);
          linebuf267 = "";
       end
    end else begin
       hitMadPrint267 = 0;
    end
  end
end


string linebuf268 = "";
logic hitMadPrint268 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc268_inst_done && ((spc268_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint268 = 1;
       linebuf268 = {linebuf268, spc268_phy_pc_w[8:1]};
       if (spc268_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 268, linebuf268);
          linebuf268 = "";
       end
    end else begin
       hitMadPrint268 = 0;
    end
  end
end


string linebuf269 = "";
logic hitMadPrint269 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc269_inst_done && ((spc269_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint269 = 1;
       linebuf269 = {linebuf269, spc269_phy_pc_w[8:1]};
       if (spc269_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 269, linebuf269);
          linebuf269 = "";
       end
    end else begin
       hitMadPrint269 = 0;
    end
  end
end


string linebuf270 = "";
logic hitMadPrint270 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc270_inst_done && ((spc270_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint270 = 1;
       linebuf270 = {linebuf270, spc270_phy_pc_w[8:1]};
       if (spc270_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 270, linebuf270);
          linebuf270 = "";
       end
    end else begin
       hitMadPrint270 = 0;
    end
  end
end


string linebuf271 = "";
logic hitMadPrint271 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc271_inst_done && ((spc271_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint271 = 1;
       linebuf271 = {linebuf271, spc271_phy_pc_w[8:1]};
       if (spc271_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 271, linebuf271);
          linebuf271 = "";
       end
    end else begin
       hitMadPrint271 = 0;
    end
  end
end


string linebuf272 = "";
logic hitMadPrint272 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc272_inst_done && ((spc272_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint272 = 1;
       linebuf272 = {linebuf272, spc272_phy_pc_w[8:1]};
       if (spc272_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 272, linebuf272);
          linebuf272 = "";
       end
    end else begin
       hitMadPrint272 = 0;
    end
  end
end


string linebuf273 = "";
logic hitMadPrint273 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc273_inst_done && ((spc273_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint273 = 1;
       linebuf273 = {linebuf273, spc273_phy_pc_w[8:1]};
       if (spc273_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 273, linebuf273);
          linebuf273 = "";
       end
    end else begin
       hitMadPrint273 = 0;
    end
  end
end


string linebuf274 = "";
logic hitMadPrint274 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc274_inst_done && ((spc274_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint274 = 1;
       linebuf274 = {linebuf274, spc274_phy_pc_w[8:1]};
       if (spc274_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 274, linebuf274);
          linebuf274 = "";
       end
    end else begin
       hitMadPrint274 = 0;
    end
  end
end


string linebuf275 = "";
logic hitMadPrint275 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc275_inst_done && ((spc275_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint275 = 1;
       linebuf275 = {linebuf275, spc275_phy_pc_w[8:1]};
       if (spc275_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 275, linebuf275);
          linebuf275 = "";
       end
    end else begin
       hitMadPrint275 = 0;
    end
  end
end


string linebuf276 = "";
logic hitMadPrint276 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc276_inst_done && ((spc276_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint276 = 1;
       linebuf276 = {linebuf276, spc276_phy_pc_w[8:1]};
       if (spc276_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 276, linebuf276);
          linebuf276 = "";
       end
    end else begin
       hitMadPrint276 = 0;
    end
  end
end


string linebuf277 = "";
logic hitMadPrint277 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc277_inst_done && ((spc277_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint277 = 1;
       linebuf277 = {linebuf277, spc277_phy_pc_w[8:1]};
       if (spc277_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 277, linebuf277);
          linebuf277 = "";
       end
    end else begin
       hitMadPrint277 = 0;
    end
  end
end


string linebuf278 = "";
logic hitMadPrint278 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc278_inst_done && ((spc278_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint278 = 1;
       linebuf278 = {linebuf278, spc278_phy_pc_w[8:1]};
       if (spc278_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 278, linebuf278);
          linebuf278 = "";
       end
    end else begin
       hitMadPrint278 = 0;
    end
  end
end


string linebuf279 = "";
logic hitMadPrint279 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc279_inst_done && ((spc279_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint279 = 1;
       linebuf279 = {linebuf279, spc279_phy_pc_w[8:1]};
       if (spc279_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 279, linebuf279);
          linebuf279 = "";
       end
    end else begin
       hitMadPrint279 = 0;
    end
  end
end


string linebuf280 = "";
logic hitMadPrint280 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc280_inst_done && ((spc280_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint280 = 1;
       linebuf280 = {linebuf280, spc280_phy_pc_w[8:1]};
       if (spc280_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 280, linebuf280);
          linebuf280 = "";
       end
    end else begin
       hitMadPrint280 = 0;
    end
  end
end


string linebuf281 = "";
logic hitMadPrint281 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc281_inst_done && ((spc281_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint281 = 1;
       linebuf281 = {linebuf281, spc281_phy_pc_w[8:1]};
       if (spc281_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 281, linebuf281);
          linebuf281 = "";
       end
    end else begin
       hitMadPrint281 = 0;
    end
  end
end


string linebuf282 = "";
logic hitMadPrint282 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc282_inst_done && ((spc282_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint282 = 1;
       linebuf282 = {linebuf282, spc282_phy_pc_w[8:1]};
       if (spc282_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 282, linebuf282);
          linebuf282 = "";
       end
    end else begin
       hitMadPrint282 = 0;
    end
  end
end


string linebuf283 = "";
logic hitMadPrint283 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc283_inst_done && ((spc283_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint283 = 1;
       linebuf283 = {linebuf283, spc283_phy_pc_w[8:1]};
       if (spc283_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 283, linebuf283);
          linebuf283 = "";
       end
    end else begin
       hitMadPrint283 = 0;
    end
  end
end


string linebuf284 = "";
logic hitMadPrint284 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc284_inst_done && ((spc284_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint284 = 1;
       linebuf284 = {linebuf284, spc284_phy_pc_w[8:1]};
       if (spc284_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 284, linebuf284);
          linebuf284 = "";
       end
    end else begin
       hitMadPrint284 = 0;
    end
  end
end


string linebuf285 = "";
logic hitMadPrint285 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc285_inst_done && ((spc285_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint285 = 1;
       linebuf285 = {linebuf285, spc285_phy_pc_w[8:1]};
       if (spc285_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 285, linebuf285);
          linebuf285 = "";
       end
    end else begin
       hitMadPrint285 = 0;
    end
  end
end


string linebuf286 = "";
logic hitMadPrint286 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc286_inst_done && ((spc286_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint286 = 1;
       linebuf286 = {linebuf286, spc286_phy_pc_w[8:1]};
       if (spc286_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 286, linebuf286);
          linebuf286 = "";
       end
    end else begin
       hitMadPrint286 = 0;
    end
  end
end


string linebuf287 = "";
logic hitMadPrint287 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc287_inst_done && ((spc287_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint287 = 1;
       linebuf287 = {linebuf287, spc287_phy_pc_w[8:1]};
       if (spc287_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 287, linebuf287);
          linebuf287 = "";
       end
    end else begin
       hitMadPrint287 = 0;
    end
  end
end


string linebuf288 = "";
logic hitMadPrint288 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc288_inst_done && ((spc288_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint288 = 1;
       linebuf288 = {linebuf288, spc288_phy_pc_w[8:1]};
       if (spc288_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 288, linebuf288);
          linebuf288 = "";
       end
    end else begin
       hitMadPrint288 = 0;
    end
  end
end


string linebuf289 = "";
logic hitMadPrint289 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc289_inst_done && ((spc289_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint289 = 1;
       linebuf289 = {linebuf289, spc289_phy_pc_w[8:1]};
       if (spc289_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 289, linebuf289);
          linebuf289 = "";
       end
    end else begin
       hitMadPrint289 = 0;
    end
  end
end


string linebuf290 = "";
logic hitMadPrint290 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc290_inst_done && ((spc290_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint290 = 1;
       linebuf290 = {linebuf290, spc290_phy_pc_w[8:1]};
       if (spc290_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 290, linebuf290);
          linebuf290 = "";
       end
    end else begin
       hitMadPrint290 = 0;
    end
  end
end


string linebuf291 = "";
logic hitMadPrint291 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc291_inst_done && ((spc291_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint291 = 1;
       linebuf291 = {linebuf291, spc291_phy_pc_w[8:1]};
       if (spc291_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 291, linebuf291);
          linebuf291 = "";
       end
    end else begin
       hitMadPrint291 = 0;
    end
  end
end


string linebuf292 = "";
logic hitMadPrint292 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc292_inst_done && ((spc292_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint292 = 1;
       linebuf292 = {linebuf292, spc292_phy_pc_w[8:1]};
       if (spc292_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 292, linebuf292);
          linebuf292 = "";
       end
    end else begin
       hitMadPrint292 = 0;
    end
  end
end


string linebuf293 = "";
logic hitMadPrint293 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc293_inst_done && ((spc293_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint293 = 1;
       linebuf293 = {linebuf293, spc293_phy_pc_w[8:1]};
       if (spc293_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 293, linebuf293);
          linebuf293 = "";
       end
    end else begin
       hitMadPrint293 = 0;
    end
  end
end


string linebuf294 = "";
logic hitMadPrint294 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc294_inst_done && ((spc294_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint294 = 1;
       linebuf294 = {linebuf294, spc294_phy_pc_w[8:1]};
       if (spc294_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 294, linebuf294);
          linebuf294 = "";
       end
    end else begin
       hitMadPrint294 = 0;
    end
  end
end


string linebuf295 = "";
logic hitMadPrint295 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc295_inst_done && ((spc295_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint295 = 1;
       linebuf295 = {linebuf295, spc295_phy_pc_w[8:1]};
       if (spc295_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 295, linebuf295);
          linebuf295 = "";
       end
    end else begin
       hitMadPrint295 = 0;
    end
  end
end


string linebuf296 = "";
logic hitMadPrint296 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc296_inst_done && ((spc296_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint296 = 1;
       linebuf296 = {linebuf296, spc296_phy_pc_w[8:1]};
       if (spc296_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 296, linebuf296);
          linebuf296 = "";
       end
    end else begin
       hitMadPrint296 = 0;
    end
  end
end


string linebuf297 = "";
logic hitMadPrint297 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc297_inst_done && ((spc297_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint297 = 1;
       linebuf297 = {linebuf297, spc297_phy_pc_w[8:1]};
       if (spc297_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 297, linebuf297);
          linebuf297 = "";
       end
    end else begin
       hitMadPrint297 = 0;
    end
  end
end


string linebuf298 = "";
logic hitMadPrint298 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc298_inst_done && ((spc298_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint298 = 1;
       linebuf298 = {linebuf298, spc298_phy_pc_w[8:1]};
       if (spc298_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 298, linebuf298);
          linebuf298 = "";
       end
    end else begin
       hitMadPrint298 = 0;
    end
  end
end


string linebuf299 = "";
logic hitMadPrint299 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc299_inst_done && ((spc299_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint299 = 1;
       linebuf299 = {linebuf299, spc299_phy_pc_w[8:1]};
       if (spc299_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 299, linebuf299);
          linebuf299 = "";
       end
    end else begin
       hitMadPrint299 = 0;
    end
  end
end


string linebuf300 = "";
logic hitMadPrint300 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc300_inst_done && ((spc300_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint300 = 1;
       linebuf300 = {linebuf300, spc300_phy_pc_w[8:1]};
       if (spc300_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 300, linebuf300);
          linebuf300 = "";
       end
    end else begin
       hitMadPrint300 = 0;
    end
  end
end


string linebuf301 = "";
logic hitMadPrint301 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc301_inst_done && ((spc301_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint301 = 1;
       linebuf301 = {linebuf301, spc301_phy_pc_w[8:1]};
       if (spc301_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 301, linebuf301);
          linebuf301 = "";
       end
    end else begin
       hitMadPrint301 = 0;
    end
  end
end


string linebuf302 = "";
logic hitMadPrint302 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc302_inst_done && ((spc302_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint302 = 1;
       linebuf302 = {linebuf302, spc302_phy_pc_w[8:1]};
       if (spc302_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 302, linebuf302);
          linebuf302 = "";
       end
    end else begin
       hitMadPrint302 = 0;
    end
  end
end


string linebuf303 = "";
logic hitMadPrint303 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc303_inst_done && ((spc303_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint303 = 1;
       linebuf303 = {linebuf303, spc303_phy_pc_w[8:1]};
       if (spc303_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 303, linebuf303);
          linebuf303 = "";
       end
    end else begin
       hitMadPrint303 = 0;
    end
  end
end


string linebuf304 = "";
logic hitMadPrint304 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc304_inst_done && ((spc304_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint304 = 1;
       linebuf304 = {linebuf304, spc304_phy_pc_w[8:1]};
       if (spc304_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 304, linebuf304);
          linebuf304 = "";
       end
    end else begin
       hitMadPrint304 = 0;
    end
  end
end


string linebuf305 = "";
logic hitMadPrint305 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc305_inst_done && ((spc305_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint305 = 1;
       linebuf305 = {linebuf305, spc305_phy_pc_w[8:1]};
       if (spc305_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 305, linebuf305);
          linebuf305 = "";
       end
    end else begin
       hitMadPrint305 = 0;
    end
  end
end


string linebuf306 = "";
logic hitMadPrint306 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc306_inst_done && ((spc306_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint306 = 1;
       linebuf306 = {linebuf306, spc306_phy_pc_w[8:1]};
       if (spc306_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 306, linebuf306);
          linebuf306 = "";
       end
    end else begin
       hitMadPrint306 = 0;
    end
  end
end


string linebuf307 = "";
logic hitMadPrint307 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc307_inst_done && ((spc307_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint307 = 1;
       linebuf307 = {linebuf307, spc307_phy_pc_w[8:1]};
       if (spc307_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 307, linebuf307);
          linebuf307 = "";
       end
    end else begin
       hitMadPrint307 = 0;
    end
  end
end


string linebuf308 = "";
logic hitMadPrint308 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc308_inst_done && ((spc308_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint308 = 1;
       linebuf308 = {linebuf308, spc308_phy_pc_w[8:1]};
       if (spc308_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 308, linebuf308);
          linebuf308 = "";
       end
    end else begin
       hitMadPrint308 = 0;
    end
  end
end


string linebuf309 = "";
logic hitMadPrint309 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc309_inst_done && ((spc309_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint309 = 1;
       linebuf309 = {linebuf309, spc309_phy_pc_w[8:1]};
       if (spc309_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 309, linebuf309);
          linebuf309 = "";
       end
    end else begin
       hitMadPrint309 = 0;
    end
  end
end


string linebuf310 = "";
logic hitMadPrint310 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc310_inst_done && ((spc310_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint310 = 1;
       linebuf310 = {linebuf310, spc310_phy_pc_w[8:1]};
       if (spc310_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 310, linebuf310);
          linebuf310 = "";
       end
    end else begin
       hitMadPrint310 = 0;
    end
  end
end


string linebuf311 = "";
logic hitMadPrint311 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc311_inst_done && ((spc311_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint311 = 1;
       linebuf311 = {linebuf311, spc311_phy_pc_w[8:1]};
       if (spc311_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 311, linebuf311);
          linebuf311 = "";
       end
    end else begin
       hitMadPrint311 = 0;
    end
  end
end


string linebuf312 = "";
logic hitMadPrint312 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc312_inst_done && ((spc312_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint312 = 1;
       linebuf312 = {linebuf312, spc312_phy_pc_w[8:1]};
       if (spc312_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 312, linebuf312);
          linebuf312 = "";
       end
    end else begin
       hitMadPrint312 = 0;
    end
  end
end


string linebuf313 = "";
logic hitMadPrint313 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc313_inst_done && ((spc313_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint313 = 1;
       linebuf313 = {linebuf313, spc313_phy_pc_w[8:1]};
       if (spc313_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 313, linebuf313);
          linebuf313 = "";
       end
    end else begin
       hitMadPrint313 = 0;
    end
  end
end


string linebuf314 = "";
logic hitMadPrint314 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc314_inst_done && ((spc314_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint314 = 1;
       linebuf314 = {linebuf314, spc314_phy_pc_w[8:1]};
       if (spc314_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 314, linebuf314);
          linebuf314 = "";
       end
    end else begin
       hitMadPrint314 = 0;
    end
  end
end


string linebuf315 = "";
logic hitMadPrint315 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc315_inst_done && ((spc315_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint315 = 1;
       linebuf315 = {linebuf315, spc315_phy_pc_w[8:1]};
       if (spc315_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 315, linebuf315);
          linebuf315 = "";
       end
    end else begin
       hitMadPrint315 = 0;
    end
  end
end


string linebuf316 = "";
logic hitMadPrint316 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc316_inst_done && ((spc316_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint316 = 1;
       linebuf316 = {linebuf316, spc316_phy_pc_w[8:1]};
       if (spc316_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 316, linebuf316);
          linebuf316 = "";
       end
    end else begin
       hitMadPrint316 = 0;
    end
  end
end


string linebuf317 = "";
logic hitMadPrint317 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc317_inst_done && ((spc317_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint317 = 1;
       linebuf317 = {linebuf317, spc317_phy_pc_w[8:1]};
       if (spc317_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 317, linebuf317);
          linebuf317 = "";
       end
    end else begin
       hitMadPrint317 = 0;
    end
  end
end


string linebuf318 = "";
logic hitMadPrint318 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc318_inst_done && ((spc318_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint318 = 1;
       linebuf318 = {linebuf318, spc318_phy_pc_w[8:1]};
       if (spc318_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 318, linebuf318);
          linebuf318 = "";
       end
    end else begin
       hitMadPrint318 = 0;
    end
  end
end


string linebuf319 = "";
logic hitMadPrint319 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc319_inst_done && ((spc319_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint319 = 1;
       linebuf319 = {linebuf319, spc319_phy_pc_w[8:1]};
       if (spc319_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 319, linebuf319);
          linebuf319 = "";
       end
    end else begin
       hitMadPrint319 = 0;
    end
  end
end


string linebuf320 = "";
logic hitMadPrint320 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc320_inst_done && ((spc320_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint320 = 1;
       linebuf320 = {linebuf320, spc320_phy_pc_w[8:1]};
       if (spc320_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 320, linebuf320);
          linebuf320 = "";
       end
    end else begin
       hitMadPrint320 = 0;
    end
  end
end


string linebuf321 = "";
logic hitMadPrint321 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc321_inst_done && ((spc321_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint321 = 1;
       linebuf321 = {linebuf321, spc321_phy_pc_w[8:1]};
       if (spc321_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 321, linebuf321);
          linebuf321 = "";
       end
    end else begin
       hitMadPrint321 = 0;
    end
  end
end


string linebuf322 = "";
logic hitMadPrint322 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc322_inst_done && ((spc322_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint322 = 1;
       linebuf322 = {linebuf322, spc322_phy_pc_w[8:1]};
       if (spc322_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 322, linebuf322);
          linebuf322 = "";
       end
    end else begin
       hitMadPrint322 = 0;
    end
  end
end


string linebuf323 = "";
logic hitMadPrint323 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc323_inst_done && ((spc323_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint323 = 1;
       linebuf323 = {linebuf323, spc323_phy_pc_w[8:1]};
       if (spc323_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 323, linebuf323);
          linebuf323 = "";
       end
    end else begin
       hitMadPrint323 = 0;
    end
  end
end


string linebuf324 = "";
logic hitMadPrint324 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc324_inst_done && ((spc324_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint324 = 1;
       linebuf324 = {linebuf324, spc324_phy_pc_w[8:1]};
       if (spc324_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 324, linebuf324);
          linebuf324 = "";
       end
    end else begin
       hitMadPrint324 = 0;
    end
  end
end


string linebuf325 = "";
logic hitMadPrint325 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc325_inst_done && ((spc325_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint325 = 1;
       linebuf325 = {linebuf325, spc325_phy_pc_w[8:1]};
       if (spc325_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 325, linebuf325);
          linebuf325 = "";
       end
    end else begin
       hitMadPrint325 = 0;
    end
  end
end


string linebuf326 = "";
logic hitMadPrint326 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc326_inst_done && ((spc326_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint326 = 1;
       linebuf326 = {linebuf326, spc326_phy_pc_w[8:1]};
       if (spc326_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 326, linebuf326);
          linebuf326 = "";
       end
    end else begin
       hitMadPrint326 = 0;
    end
  end
end


string linebuf327 = "";
logic hitMadPrint327 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc327_inst_done && ((spc327_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint327 = 1;
       linebuf327 = {linebuf327, spc327_phy_pc_w[8:1]};
       if (spc327_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 327, linebuf327);
          linebuf327 = "";
       end
    end else begin
       hitMadPrint327 = 0;
    end
  end
end


string linebuf328 = "";
logic hitMadPrint328 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc328_inst_done && ((spc328_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint328 = 1;
       linebuf328 = {linebuf328, spc328_phy_pc_w[8:1]};
       if (spc328_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 328, linebuf328);
          linebuf328 = "";
       end
    end else begin
       hitMadPrint328 = 0;
    end
  end
end


string linebuf329 = "";
logic hitMadPrint329 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc329_inst_done && ((spc329_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint329 = 1;
       linebuf329 = {linebuf329, spc329_phy_pc_w[8:1]};
       if (spc329_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 329, linebuf329);
          linebuf329 = "";
       end
    end else begin
       hitMadPrint329 = 0;
    end
  end
end


string linebuf330 = "";
logic hitMadPrint330 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc330_inst_done && ((spc330_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint330 = 1;
       linebuf330 = {linebuf330, spc330_phy_pc_w[8:1]};
       if (spc330_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 330, linebuf330);
          linebuf330 = "";
       end
    end else begin
       hitMadPrint330 = 0;
    end
  end
end


string linebuf331 = "";
logic hitMadPrint331 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc331_inst_done && ((spc331_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint331 = 1;
       linebuf331 = {linebuf331, spc331_phy_pc_w[8:1]};
       if (spc331_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 331, linebuf331);
          linebuf331 = "";
       end
    end else begin
       hitMadPrint331 = 0;
    end
  end
end


string linebuf332 = "";
logic hitMadPrint332 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc332_inst_done && ((spc332_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint332 = 1;
       linebuf332 = {linebuf332, spc332_phy_pc_w[8:1]};
       if (spc332_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 332, linebuf332);
          linebuf332 = "";
       end
    end else begin
       hitMadPrint332 = 0;
    end
  end
end


string linebuf333 = "";
logic hitMadPrint333 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc333_inst_done && ((spc333_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint333 = 1;
       linebuf333 = {linebuf333, spc333_phy_pc_w[8:1]};
       if (spc333_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 333, linebuf333);
          linebuf333 = "";
       end
    end else begin
       hitMadPrint333 = 0;
    end
  end
end


string linebuf334 = "";
logic hitMadPrint334 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc334_inst_done && ((spc334_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint334 = 1;
       linebuf334 = {linebuf334, spc334_phy_pc_w[8:1]};
       if (spc334_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 334, linebuf334);
          linebuf334 = "";
       end
    end else begin
       hitMadPrint334 = 0;
    end
  end
end


string linebuf335 = "";
logic hitMadPrint335 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc335_inst_done && ((spc335_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint335 = 1;
       linebuf335 = {linebuf335, spc335_phy_pc_w[8:1]};
       if (spc335_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 335, linebuf335);
          linebuf335 = "";
       end
    end else begin
       hitMadPrint335 = 0;
    end
  end
end


string linebuf336 = "";
logic hitMadPrint336 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc336_inst_done && ((spc336_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint336 = 1;
       linebuf336 = {linebuf336, spc336_phy_pc_w[8:1]};
       if (spc336_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 336, linebuf336);
          linebuf336 = "";
       end
    end else begin
       hitMadPrint336 = 0;
    end
  end
end


string linebuf337 = "";
logic hitMadPrint337 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc337_inst_done && ((spc337_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint337 = 1;
       linebuf337 = {linebuf337, spc337_phy_pc_w[8:1]};
       if (spc337_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 337, linebuf337);
          linebuf337 = "";
       end
    end else begin
       hitMadPrint337 = 0;
    end
  end
end


string linebuf338 = "";
logic hitMadPrint338 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc338_inst_done && ((spc338_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint338 = 1;
       linebuf338 = {linebuf338, spc338_phy_pc_w[8:1]};
       if (spc338_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 338, linebuf338);
          linebuf338 = "";
       end
    end else begin
       hitMadPrint338 = 0;
    end
  end
end


string linebuf339 = "";
logic hitMadPrint339 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc339_inst_done && ((spc339_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint339 = 1;
       linebuf339 = {linebuf339, spc339_phy_pc_w[8:1]};
       if (spc339_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 339, linebuf339);
          linebuf339 = "";
       end
    end else begin
       hitMadPrint339 = 0;
    end
  end
end


string linebuf340 = "";
logic hitMadPrint340 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc340_inst_done && ((spc340_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint340 = 1;
       linebuf340 = {linebuf340, spc340_phy_pc_w[8:1]};
       if (spc340_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 340, linebuf340);
          linebuf340 = "";
       end
    end else begin
       hitMadPrint340 = 0;
    end
  end
end


string linebuf341 = "";
logic hitMadPrint341 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc341_inst_done && ((spc341_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint341 = 1;
       linebuf341 = {linebuf341, spc341_phy_pc_w[8:1]};
       if (spc341_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 341, linebuf341);
          linebuf341 = "";
       end
    end else begin
       hitMadPrint341 = 0;
    end
  end
end


string linebuf342 = "";
logic hitMadPrint342 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc342_inst_done && ((spc342_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint342 = 1;
       linebuf342 = {linebuf342, spc342_phy_pc_w[8:1]};
       if (spc342_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 342, linebuf342);
          linebuf342 = "";
       end
    end else begin
       hitMadPrint342 = 0;
    end
  end
end


string linebuf343 = "";
logic hitMadPrint343 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc343_inst_done && ((spc343_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint343 = 1;
       linebuf343 = {linebuf343, spc343_phy_pc_w[8:1]};
       if (spc343_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 343, linebuf343);
          linebuf343 = "";
       end
    end else begin
       hitMadPrint343 = 0;
    end
  end
end


string linebuf344 = "";
logic hitMadPrint344 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc344_inst_done && ((spc344_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint344 = 1;
       linebuf344 = {linebuf344, spc344_phy_pc_w[8:1]};
       if (spc344_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 344, linebuf344);
          linebuf344 = "";
       end
    end else begin
       hitMadPrint344 = 0;
    end
  end
end


string linebuf345 = "";
logic hitMadPrint345 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc345_inst_done && ((spc345_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint345 = 1;
       linebuf345 = {linebuf345, spc345_phy_pc_w[8:1]};
       if (spc345_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 345, linebuf345);
          linebuf345 = "";
       end
    end else begin
       hitMadPrint345 = 0;
    end
  end
end


string linebuf346 = "";
logic hitMadPrint346 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc346_inst_done && ((spc346_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint346 = 1;
       linebuf346 = {linebuf346, spc346_phy_pc_w[8:1]};
       if (spc346_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 346, linebuf346);
          linebuf346 = "";
       end
    end else begin
       hitMadPrint346 = 0;
    end
  end
end


string linebuf347 = "";
logic hitMadPrint347 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc347_inst_done && ((spc347_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint347 = 1;
       linebuf347 = {linebuf347, spc347_phy_pc_w[8:1]};
       if (spc347_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 347, linebuf347);
          linebuf347 = "";
       end
    end else begin
       hitMadPrint347 = 0;
    end
  end
end


string linebuf348 = "";
logic hitMadPrint348 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc348_inst_done && ((spc348_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint348 = 1;
       linebuf348 = {linebuf348, spc348_phy_pc_w[8:1]};
       if (spc348_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 348, linebuf348);
          linebuf348 = "";
       end
    end else begin
       hitMadPrint348 = 0;
    end
  end
end


string linebuf349 = "";
logic hitMadPrint349 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc349_inst_done && ((spc349_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint349 = 1;
       linebuf349 = {linebuf349, spc349_phy_pc_w[8:1]};
       if (spc349_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 349, linebuf349);
          linebuf349 = "";
       end
    end else begin
       hitMadPrint349 = 0;
    end
  end
end


string linebuf350 = "";
logic hitMadPrint350 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc350_inst_done && ((spc350_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint350 = 1;
       linebuf350 = {linebuf350, spc350_phy_pc_w[8:1]};
       if (spc350_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 350, linebuf350);
          linebuf350 = "";
       end
    end else begin
       hitMadPrint350 = 0;
    end
  end
end


string linebuf351 = "";
logic hitMadPrint351 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc351_inst_done && ((spc351_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint351 = 1;
       linebuf351 = {linebuf351, spc351_phy_pc_w[8:1]};
       if (spc351_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 351, linebuf351);
          linebuf351 = "";
       end
    end else begin
       hitMadPrint351 = 0;
    end
  end
end


string linebuf352 = "";
logic hitMadPrint352 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc352_inst_done && ((spc352_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint352 = 1;
       linebuf352 = {linebuf352, spc352_phy_pc_w[8:1]};
       if (spc352_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 352, linebuf352);
          linebuf352 = "";
       end
    end else begin
       hitMadPrint352 = 0;
    end
  end
end


string linebuf353 = "";
logic hitMadPrint353 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc353_inst_done && ((spc353_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint353 = 1;
       linebuf353 = {linebuf353, spc353_phy_pc_w[8:1]};
       if (spc353_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 353, linebuf353);
          linebuf353 = "";
       end
    end else begin
       hitMadPrint353 = 0;
    end
  end
end


string linebuf354 = "";
logic hitMadPrint354 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc354_inst_done && ((spc354_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint354 = 1;
       linebuf354 = {linebuf354, spc354_phy_pc_w[8:1]};
       if (spc354_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 354, linebuf354);
          linebuf354 = "";
       end
    end else begin
       hitMadPrint354 = 0;
    end
  end
end


string linebuf355 = "";
logic hitMadPrint355 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc355_inst_done && ((spc355_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint355 = 1;
       linebuf355 = {linebuf355, spc355_phy_pc_w[8:1]};
       if (spc355_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 355, linebuf355);
          linebuf355 = "";
       end
    end else begin
       hitMadPrint355 = 0;
    end
  end
end


string linebuf356 = "";
logic hitMadPrint356 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc356_inst_done && ((spc356_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint356 = 1;
       linebuf356 = {linebuf356, spc356_phy_pc_w[8:1]};
       if (spc356_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 356, linebuf356);
          linebuf356 = "";
       end
    end else begin
       hitMadPrint356 = 0;
    end
  end
end


string linebuf357 = "";
logic hitMadPrint357 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc357_inst_done && ((spc357_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint357 = 1;
       linebuf357 = {linebuf357, spc357_phy_pc_w[8:1]};
       if (spc357_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 357, linebuf357);
          linebuf357 = "";
       end
    end else begin
       hitMadPrint357 = 0;
    end
  end
end


string linebuf358 = "";
logic hitMadPrint358 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc358_inst_done && ((spc358_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint358 = 1;
       linebuf358 = {linebuf358, spc358_phy_pc_w[8:1]};
       if (spc358_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 358, linebuf358);
          linebuf358 = "";
       end
    end else begin
       hitMadPrint358 = 0;
    end
  end
end


string linebuf359 = "";
logic hitMadPrint359 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc359_inst_done && ((spc359_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint359 = 1;
       linebuf359 = {linebuf359, spc359_phy_pc_w[8:1]};
       if (spc359_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 359, linebuf359);
          linebuf359 = "";
       end
    end else begin
       hitMadPrint359 = 0;
    end
  end
end


string linebuf360 = "";
logic hitMadPrint360 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc360_inst_done && ((spc360_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint360 = 1;
       linebuf360 = {linebuf360, spc360_phy_pc_w[8:1]};
       if (spc360_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 360, linebuf360);
          linebuf360 = "";
       end
    end else begin
       hitMadPrint360 = 0;
    end
  end
end


string linebuf361 = "";
logic hitMadPrint361 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc361_inst_done && ((spc361_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint361 = 1;
       linebuf361 = {linebuf361, spc361_phy_pc_w[8:1]};
       if (spc361_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 361, linebuf361);
          linebuf361 = "";
       end
    end else begin
       hitMadPrint361 = 0;
    end
  end
end


string linebuf362 = "";
logic hitMadPrint362 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc362_inst_done && ((spc362_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint362 = 1;
       linebuf362 = {linebuf362, spc362_phy_pc_w[8:1]};
       if (spc362_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 362, linebuf362);
          linebuf362 = "";
       end
    end else begin
       hitMadPrint362 = 0;
    end
  end
end


string linebuf363 = "";
logic hitMadPrint363 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc363_inst_done && ((spc363_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint363 = 1;
       linebuf363 = {linebuf363, spc363_phy_pc_w[8:1]};
       if (spc363_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 363, linebuf363);
          linebuf363 = "";
       end
    end else begin
       hitMadPrint363 = 0;
    end
  end
end


string linebuf364 = "";
logic hitMadPrint364 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc364_inst_done && ((spc364_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint364 = 1;
       linebuf364 = {linebuf364, spc364_phy_pc_w[8:1]};
       if (spc364_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 364, linebuf364);
          linebuf364 = "";
       end
    end else begin
       hitMadPrint364 = 0;
    end
  end
end


string linebuf365 = "";
logic hitMadPrint365 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc365_inst_done && ((spc365_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint365 = 1;
       linebuf365 = {linebuf365, spc365_phy_pc_w[8:1]};
       if (spc365_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 365, linebuf365);
          linebuf365 = "";
       end
    end else begin
       hitMadPrint365 = 0;
    end
  end
end


string linebuf366 = "";
logic hitMadPrint366 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc366_inst_done && ((spc366_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint366 = 1;
       linebuf366 = {linebuf366, spc366_phy_pc_w[8:1]};
       if (spc366_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 366, linebuf366);
          linebuf366 = "";
       end
    end else begin
       hitMadPrint366 = 0;
    end
  end
end


string linebuf367 = "";
logic hitMadPrint367 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc367_inst_done && ((spc367_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint367 = 1;
       linebuf367 = {linebuf367, spc367_phy_pc_w[8:1]};
       if (spc367_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 367, linebuf367);
          linebuf367 = "";
       end
    end else begin
       hitMadPrint367 = 0;
    end
  end
end


string linebuf368 = "";
logic hitMadPrint368 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc368_inst_done && ((spc368_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint368 = 1;
       linebuf368 = {linebuf368, spc368_phy_pc_w[8:1]};
       if (spc368_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 368, linebuf368);
          linebuf368 = "";
       end
    end else begin
       hitMadPrint368 = 0;
    end
  end
end


string linebuf369 = "";
logic hitMadPrint369 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc369_inst_done && ((spc369_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint369 = 1;
       linebuf369 = {linebuf369, spc369_phy_pc_w[8:1]};
       if (spc369_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 369, linebuf369);
          linebuf369 = "";
       end
    end else begin
       hitMadPrint369 = 0;
    end
  end
end


string linebuf370 = "";
logic hitMadPrint370 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc370_inst_done && ((spc370_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint370 = 1;
       linebuf370 = {linebuf370, spc370_phy_pc_w[8:1]};
       if (spc370_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 370, linebuf370);
          linebuf370 = "";
       end
    end else begin
       hitMadPrint370 = 0;
    end
  end
end


string linebuf371 = "";
logic hitMadPrint371 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc371_inst_done && ((spc371_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint371 = 1;
       linebuf371 = {linebuf371, spc371_phy_pc_w[8:1]};
       if (spc371_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 371, linebuf371);
          linebuf371 = "";
       end
    end else begin
       hitMadPrint371 = 0;
    end
  end
end


string linebuf372 = "";
logic hitMadPrint372 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc372_inst_done && ((spc372_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint372 = 1;
       linebuf372 = {linebuf372, spc372_phy_pc_w[8:1]};
       if (spc372_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 372, linebuf372);
          linebuf372 = "";
       end
    end else begin
       hitMadPrint372 = 0;
    end
  end
end


string linebuf373 = "";
logic hitMadPrint373 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc373_inst_done && ((spc373_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint373 = 1;
       linebuf373 = {linebuf373, spc373_phy_pc_w[8:1]};
       if (spc373_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 373, linebuf373);
          linebuf373 = "";
       end
    end else begin
       hitMadPrint373 = 0;
    end
  end
end


string linebuf374 = "";
logic hitMadPrint374 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc374_inst_done && ((spc374_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint374 = 1;
       linebuf374 = {linebuf374, spc374_phy_pc_w[8:1]};
       if (spc374_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 374, linebuf374);
          linebuf374 = "";
       end
    end else begin
       hitMadPrint374 = 0;
    end
  end
end


string linebuf375 = "";
logic hitMadPrint375 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc375_inst_done && ((spc375_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint375 = 1;
       linebuf375 = {linebuf375, spc375_phy_pc_w[8:1]};
       if (spc375_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 375, linebuf375);
          linebuf375 = "";
       end
    end else begin
       hitMadPrint375 = 0;
    end
  end
end


string linebuf376 = "";
logic hitMadPrint376 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc376_inst_done && ((spc376_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint376 = 1;
       linebuf376 = {linebuf376, spc376_phy_pc_w[8:1]};
       if (spc376_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 376, linebuf376);
          linebuf376 = "";
       end
    end else begin
       hitMadPrint376 = 0;
    end
  end
end


string linebuf377 = "";
logic hitMadPrint377 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc377_inst_done && ((spc377_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint377 = 1;
       linebuf377 = {linebuf377, spc377_phy_pc_w[8:1]};
       if (spc377_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 377, linebuf377);
          linebuf377 = "";
       end
    end else begin
       hitMadPrint377 = 0;
    end
  end
end


string linebuf378 = "";
logic hitMadPrint378 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc378_inst_done && ((spc378_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint378 = 1;
       linebuf378 = {linebuf378, spc378_phy_pc_w[8:1]};
       if (spc378_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 378, linebuf378);
          linebuf378 = "";
       end
    end else begin
       hitMadPrint378 = 0;
    end
  end
end


string linebuf379 = "";
logic hitMadPrint379 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc379_inst_done && ((spc379_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint379 = 1;
       linebuf379 = {linebuf379, spc379_phy_pc_w[8:1]};
       if (spc379_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 379, linebuf379);
          linebuf379 = "";
       end
    end else begin
       hitMadPrint379 = 0;
    end
  end
end


string linebuf380 = "";
logic hitMadPrint380 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc380_inst_done && ((spc380_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint380 = 1;
       linebuf380 = {linebuf380, spc380_phy_pc_w[8:1]};
       if (spc380_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 380, linebuf380);
          linebuf380 = "";
       end
    end else begin
       hitMadPrint380 = 0;
    end
  end
end


string linebuf381 = "";
logic hitMadPrint381 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc381_inst_done && ((spc381_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint381 = 1;
       linebuf381 = {linebuf381, spc381_phy_pc_w[8:1]};
       if (spc381_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 381, linebuf381);
          linebuf381 = "";
       end
    end else begin
       hitMadPrint381 = 0;
    end
  end
end


string linebuf382 = "";
logic hitMadPrint382 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc382_inst_done && ((spc382_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint382 = 1;
       linebuf382 = {linebuf382, spc382_phy_pc_w[8:1]};
       if (spc382_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 382, linebuf382);
          linebuf382 = "";
       end
    end else begin
       hitMadPrint382 = 0;
    end
  end
end


string linebuf383 = "";
logic hitMadPrint383 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc383_inst_done && ((spc383_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint383 = 1;
       linebuf383 = {linebuf383, spc383_phy_pc_w[8:1]};
       if (spc383_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 383, linebuf383);
          linebuf383 = "";
       end
    end else begin
       hitMadPrint383 = 0;
    end
  end
end


string linebuf384 = "";
logic hitMadPrint384 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc384_inst_done && ((spc384_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint384 = 1;
       linebuf384 = {linebuf384, spc384_phy_pc_w[8:1]};
       if (spc384_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 384, linebuf384);
          linebuf384 = "";
       end
    end else begin
       hitMadPrint384 = 0;
    end
  end
end


string linebuf385 = "";
logic hitMadPrint385 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc385_inst_done && ((spc385_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint385 = 1;
       linebuf385 = {linebuf385, spc385_phy_pc_w[8:1]};
       if (spc385_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 385, linebuf385);
          linebuf385 = "";
       end
    end else begin
       hitMadPrint385 = 0;
    end
  end
end


string linebuf386 = "";
logic hitMadPrint386 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc386_inst_done && ((spc386_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint386 = 1;
       linebuf386 = {linebuf386, spc386_phy_pc_w[8:1]};
       if (spc386_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 386, linebuf386);
          linebuf386 = "";
       end
    end else begin
       hitMadPrint386 = 0;
    end
  end
end


string linebuf387 = "";
logic hitMadPrint387 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc387_inst_done && ((spc387_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint387 = 1;
       linebuf387 = {linebuf387, spc387_phy_pc_w[8:1]};
       if (spc387_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 387, linebuf387);
          linebuf387 = "";
       end
    end else begin
       hitMadPrint387 = 0;
    end
  end
end


string linebuf388 = "";
logic hitMadPrint388 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc388_inst_done && ((spc388_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint388 = 1;
       linebuf388 = {linebuf388, spc388_phy_pc_w[8:1]};
       if (spc388_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 388, linebuf388);
          linebuf388 = "";
       end
    end else begin
       hitMadPrint388 = 0;
    end
  end
end


string linebuf389 = "";
logic hitMadPrint389 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc389_inst_done && ((spc389_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint389 = 1;
       linebuf389 = {linebuf389, spc389_phy_pc_w[8:1]};
       if (spc389_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 389, linebuf389);
          linebuf389 = "";
       end
    end else begin
       hitMadPrint389 = 0;
    end
  end
end


string linebuf390 = "";
logic hitMadPrint390 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc390_inst_done && ((spc390_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint390 = 1;
       linebuf390 = {linebuf390, spc390_phy_pc_w[8:1]};
       if (spc390_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 390, linebuf390);
          linebuf390 = "";
       end
    end else begin
       hitMadPrint390 = 0;
    end
  end
end


string linebuf391 = "";
logic hitMadPrint391 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc391_inst_done && ((spc391_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint391 = 1;
       linebuf391 = {linebuf391, spc391_phy_pc_w[8:1]};
       if (spc391_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 391, linebuf391);
          linebuf391 = "";
       end
    end else begin
       hitMadPrint391 = 0;
    end
  end
end


string linebuf392 = "";
logic hitMadPrint392 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc392_inst_done && ((spc392_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint392 = 1;
       linebuf392 = {linebuf392, spc392_phy_pc_w[8:1]};
       if (spc392_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 392, linebuf392);
          linebuf392 = "";
       end
    end else begin
       hitMadPrint392 = 0;
    end
  end
end


string linebuf393 = "";
logic hitMadPrint393 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc393_inst_done && ((spc393_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint393 = 1;
       linebuf393 = {linebuf393, spc393_phy_pc_w[8:1]};
       if (spc393_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 393, linebuf393);
          linebuf393 = "";
       end
    end else begin
       hitMadPrint393 = 0;
    end
  end
end


string linebuf394 = "";
logic hitMadPrint394 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc394_inst_done && ((spc394_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint394 = 1;
       linebuf394 = {linebuf394, spc394_phy_pc_w[8:1]};
       if (spc394_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 394, linebuf394);
          linebuf394 = "";
       end
    end else begin
       hitMadPrint394 = 0;
    end
  end
end


string linebuf395 = "";
logic hitMadPrint395 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc395_inst_done && ((spc395_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint395 = 1;
       linebuf395 = {linebuf395, spc395_phy_pc_w[8:1]};
       if (spc395_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 395, linebuf395);
          linebuf395 = "";
       end
    end else begin
       hitMadPrint395 = 0;
    end
  end
end


string linebuf396 = "";
logic hitMadPrint396 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc396_inst_done && ((spc396_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint396 = 1;
       linebuf396 = {linebuf396, spc396_phy_pc_w[8:1]};
       if (spc396_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 396, linebuf396);
          linebuf396 = "";
       end
    end else begin
       hitMadPrint396 = 0;
    end
  end
end


string linebuf397 = "";
logic hitMadPrint397 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc397_inst_done && ((spc397_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint397 = 1;
       linebuf397 = {linebuf397, spc397_phy_pc_w[8:1]};
       if (spc397_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 397, linebuf397);
          linebuf397 = "";
       end
    end else begin
       hitMadPrint397 = 0;
    end
  end
end


string linebuf398 = "";
logic hitMadPrint398 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc398_inst_done && ((spc398_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint398 = 1;
       linebuf398 = {linebuf398, spc398_phy_pc_w[8:1]};
       if (spc398_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 398, linebuf398);
          linebuf398 = "";
       end
    end else begin
       hitMadPrint398 = 0;
    end
  end
end


string linebuf399 = "";
logic hitMadPrint399 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc399_inst_done && ((spc399_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint399 = 1;
       linebuf399 = {linebuf399, spc399_phy_pc_w[8:1]};
       if (spc399_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 399, linebuf399);
          linebuf399 = "";
       end
    end else begin
       hitMadPrint399 = 0;
    end
  end
end


string linebuf400 = "";
logic hitMadPrint400 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc400_inst_done && ((spc400_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint400 = 1;
       linebuf400 = {linebuf400, spc400_phy_pc_w[8:1]};
       if (spc400_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 400, linebuf400);
          linebuf400 = "";
       end
    end else begin
       hitMadPrint400 = 0;
    end
  end
end


string linebuf401 = "";
logic hitMadPrint401 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc401_inst_done && ((spc401_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint401 = 1;
       linebuf401 = {linebuf401, spc401_phy_pc_w[8:1]};
       if (spc401_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 401, linebuf401);
          linebuf401 = "";
       end
    end else begin
       hitMadPrint401 = 0;
    end
  end
end


string linebuf402 = "";
logic hitMadPrint402 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc402_inst_done && ((spc402_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint402 = 1;
       linebuf402 = {linebuf402, spc402_phy_pc_w[8:1]};
       if (spc402_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 402, linebuf402);
          linebuf402 = "";
       end
    end else begin
       hitMadPrint402 = 0;
    end
  end
end


string linebuf403 = "";
logic hitMadPrint403 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc403_inst_done && ((spc403_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint403 = 1;
       linebuf403 = {linebuf403, spc403_phy_pc_w[8:1]};
       if (spc403_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 403, linebuf403);
          linebuf403 = "";
       end
    end else begin
       hitMadPrint403 = 0;
    end
  end
end


string linebuf404 = "";
logic hitMadPrint404 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc404_inst_done && ((spc404_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint404 = 1;
       linebuf404 = {linebuf404, spc404_phy_pc_w[8:1]};
       if (spc404_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 404, linebuf404);
          linebuf404 = "";
       end
    end else begin
       hitMadPrint404 = 0;
    end
  end
end


string linebuf405 = "";
logic hitMadPrint405 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc405_inst_done && ((spc405_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint405 = 1;
       linebuf405 = {linebuf405, spc405_phy_pc_w[8:1]};
       if (spc405_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 405, linebuf405);
          linebuf405 = "";
       end
    end else begin
       hitMadPrint405 = 0;
    end
  end
end


string linebuf406 = "";
logic hitMadPrint406 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc406_inst_done && ((spc406_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint406 = 1;
       linebuf406 = {linebuf406, spc406_phy_pc_w[8:1]};
       if (spc406_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 406, linebuf406);
          linebuf406 = "";
       end
    end else begin
       hitMadPrint406 = 0;
    end
  end
end


string linebuf407 = "";
logic hitMadPrint407 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc407_inst_done && ((spc407_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint407 = 1;
       linebuf407 = {linebuf407, spc407_phy_pc_w[8:1]};
       if (spc407_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 407, linebuf407);
          linebuf407 = "";
       end
    end else begin
       hitMadPrint407 = 0;
    end
  end
end


string linebuf408 = "";
logic hitMadPrint408 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc408_inst_done && ((spc408_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint408 = 1;
       linebuf408 = {linebuf408, spc408_phy_pc_w[8:1]};
       if (spc408_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 408, linebuf408);
          linebuf408 = "";
       end
    end else begin
       hitMadPrint408 = 0;
    end
  end
end


string linebuf409 = "";
logic hitMadPrint409 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc409_inst_done && ((spc409_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint409 = 1;
       linebuf409 = {linebuf409, spc409_phy_pc_w[8:1]};
       if (spc409_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 409, linebuf409);
          linebuf409 = "";
       end
    end else begin
       hitMadPrint409 = 0;
    end
  end
end


string linebuf410 = "";
logic hitMadPrint410 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc410_inst_done && ((spc410_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint410 = 1;
       linebuf410 = {linebuf410, spc410_phy_pc_w[8:1]};
       if (spc410_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 410, linebuf410);
          linebuf410 = "";
       end
    end else begin
       hitMadPrint410 = 0;
    end
  end
end


string linebuf411 = "";
logic hitMadPrint411 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc411_inst_done && ((spc411_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint411 = 1;
       linebuf411 = {linebuf411, spc411_phy_pc_w[8:1]};
       if (spc411_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 411, linebuf411);
          linebuf411 = "";
       end
    end else begin
       hitMadPrint411 = 0;
    end
  end
end


string linebuf412 = "";
logic hitMadPrint412 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc412_inst_done && ((spc412_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint412 = 1;
       linebuf412 = {linebuf412, spc412_phy_pc_w[8:1]};
       if (spc412_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 412, linebuf412);
          linebuf412 = "";
       end
    end else begin
       hitMadPrint412 = 0;
    end
  end
end


string linebuf413 = "";
logic hitMadPrint413 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc413_inst_done && ((spc413_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint413 = 1;
       linebuf413 = {linebuf413, spc413_phy_pc_w[8:1]};
       if (spc413_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 413, linebuf413);
          linebuf413 = "";
       end
    end else begin
       hitMadPrint413 = 0;
    end
  end
end


string linebuf414 = "";
logic hitMadPrint414 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc414_inst_done && ((spc414_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint414 = 1;
       linebuf414 = {linebuf414, spc414_phy_pc_w[8:1]};
       if (spc414_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 414, linebuf414);
          linebuf414 = "";
       end
    end else begin
       hitMadPrint414 = 0;
    end
  end
end


string linebuf415 = "";
logic hitMadPrint415 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc415_inst_done && ((spc415_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint415 = 1;
       linebuf415 = {linebuf415, spc415_phy_pc_w[8:1]};
       if (spc415_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 415, linebuf415);
          linebuf415 = "";
       end
    end else begin
       hitMadPrint415 = 0;
    end
  end
end


string linebuf416 = "";
logic hitMadPrint416 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc416_inst_done && ((spc416_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint416 = 1;
       linebuf416 = {linebuf416, spc416_phy_pc_w[8:1]};
       if (spc416_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 416, linebuf416);
          linebuf416 = "";
       end
    end else begin
       hitMadPrint416 = 0;
    end
  end
end


string linebuf417 = "";
logic hitMadPrint417 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc417_inst_done && ((spc417_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint417 = 1;
       linebuf417 = {linebuf417, spc417_phy_pc_w[8:1]};
       if (spc417_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 417, linebuf417);
          linebuf417 = "";
       end
    end else begin
       hitMadPrint417 = 0;
    end
  end
end


string linebuf418 = "";
logic hitMadPrint418 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc418_inst_done && ((spc418_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint418 = 1;
       linebuf418 = {linebuf418, spc418_phy_pc_w[8:1]};
       if (spc418_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 418, linebuf418);
          linebuf418 = "";
       end
    end else begin
       hitMadPrint418 = 0;
    end
  end
end


string linebuf419 = "";
logic hitMadPrint419 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc419_inst_done && ((spc419_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint419 = 1;
       linebuf419 = {linebuf419, spc419_phy_pc_w[8:1]};
       if (spc419_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 419, linebuf419);
          linebuf419 = "";
       end
    end else begin
       hitMadPrint419 = 0;
    end
  end
end


string linebuf420 = "";
logic hitMadPrint420 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc420_inst_done && ((spc420_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint420 = 1;
       linebuf420 = {linebuf420, spc420_phy_pc_w[8:1]};
       if (spc420_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 420, linebuf420);
          linebuf420 = "";
       end
    end else begin
       hitMadPrint420 = 0;
    end
  end
end


string linebuf421 = "";
logic hitMadPrint421 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc421_inst_done && ((spc421_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint421 = 1;
       linebuf421 = {linebuf421, spc421_phy_pc_w[8:1]};
       if (spc421_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 421, linebuf421);
          linebuf421 = "";
       end
    end else begin
       hitMadPrint421 = 0;
    end
  end
end


string linebuf422 = "";
logic hitMadPrint422 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc422_inst_done && ((spc422_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint422 = 1;
       linebuf422 = {linebuf422, spc422_phy_pc_w[8:1]};
       if (spc422_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 422, linebuf422);
          linebuf422 = "";
       end
    end else begin
       hitMadPrint422 = 0;
    end
  end
end


string linebuf423 = "";
logic hitMadPrint423 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc423_inst_done && ((spc423_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint423 = 1;
       linebuf423 = {linebuf423, spc423_phy_pc_w[8:1]};
       if (spc423_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 423, linebuf423);
          linebuf423 = "";
       end
    end else begin
       hitMadPrint423 = 0;
    end
  end
end


string linebuf424 = "";
logic hitMadPrint424 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc424_inst_done && ((spc424_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint424 = 1;
       linebuf424 = {linebuf424, spc424_phy_pc_w[8:1]};
       if (spc424_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 424, linebuf424);
          linebuf424 = "";
       end
    end else begin
       hitMadPrint424 = 0;
    end
  end
end


string linebuf425 = "";
logic hitMadPrint425 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc425_inst_done && ((spc425_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint425 = 1;
       linebuf425 = {linebuf425, spc425_phy_pc_w[8:1]};
       if (spc425_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 425, linebuf425);
          linebuf425 = "";
       end
    end else begin
       hitMadPrint425 = 0;
    end
  end
end


string linebuf426 = "";
logic hitMadPrint426 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc426_inst_done && ((spc426_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint426 = 1;
       linebuf426 = {linebuf426, spc426_phy_pc_w[8:1]};
       if (spc426_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 426, linebuf426);
          linebuf426 = "";
       end
    end else begin
       hitMadPrint426 = 0;
    end
  end
end


string linebuf427 = "";
logic hitMadPrint427 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc427_inst_done && ((spc427_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint427 = 1;
       linebuf427 = {linebuf427, spc427_phy_pc_w[8:1]};
       if (spc427_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 427, linebuf427);
          linebuf427 = "";
       end
    end else begin
       hitMadPrint427 = 0;
    end
  end
end


string linebuf428 = "";
logic hitMadPrint428 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc428_inst_done && ((spc428_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint428 = 1;
       linebuf428 = {linebuf428, spc428_phy_pc_w[8:1]};
       if (spc428_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 428, linebuf428);
          linebuf428 = "";
       end
    end else begin
       hitMadPrint428 = 0;
    end
  end
end


string linebuf429 = "";
logic hitMadPrint429 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc429_inst_done && ((spc429_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint429 = 1;
       linebuf429 = {linebuf429, spc429_phy_pc_w[8:1]};
       if (spc429_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 429, linebuf429);
          linebuf429 = "";
       end
    end else begin
       hitMadPrint429 = 0;
    end
  end
end


string linebuf430 = "";
logic hitMadPrint430 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc430_inst_done && ((spc430_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint430 = 1;
       linebuf430 = {linebuf430, spc430_phy_pc_w[8:1]};
       if (spc430_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 430, linebuf430);
          linebuf430 = "";
       end
    end else begin
       hitMadPrint430 = 0;
    end
  end
end


string linebuf431 = "";
logic hitMadPrint431 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc431_inst_done && ((spc431_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint431 = 1;
       linebuf431 = {linebuf431, spc431_phy_pc_w[8:1]};
       if (spc431_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 431, linebuf431);
          linebuf431 = "";
       end
    end else begin
       hitMadPrint431 = 0;
    end
  end
end


string linebuf432 = "";
logic hitMadPrint432 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc432_inst_done && ((spc432_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint432 = 1;
       linebuf432 = {linebuf432, spc432_phy_pc_w[8:1]};
       if (spc432_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 432, linebuf432);
          linebuf432 = "";
       end
    end else begin
       hitMadPrint432 = 0;
    end
  end
end


string linebuf433 = "";
logic hitMadPrint433 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc433_inst_done && ((spc433_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint433 = 1;
       linebuf433 = {linebuf433, spc433_phy_pc_w[8:1]};
       if (spc433_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 433, linebuf433);
          linebuf433 = "";
       end
    end else begin
       hitMadPrint433 = 0;
    end
  end
end


string linebuf434 = "";
logic hitMadPrint434 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc434_inst_done && ((spc434_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint434 = 1;
       linebuf434 = {linebuf434, spc434_phy_pc_w[8:1]};
       if (spc434_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 434, linebuf434);
          linebuf434 = "";
       end
    end else begin
       hitMadPrint434 = 0;
    end
  end
end


string linebuf435 = "";
logic hitMadPrint435 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc435_inst_done && ((spc435_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint435 = 1;
       linebuf435 = {linebuf435, spc435_phy_pc_w[8:1]};
       if (spc435_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 435, linebuf435);
          linebuf435 = "";
       end
    end else begin
       hitMadPrint435 = 0;
    end
  end
end


string linebuf436 = "";
logic hitMadPrint436 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc436_inst_done && ((spc436_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint436 = 1;
       linebuf436 = {linebuf436, spc436_phy_pc_w[8:1]};
       if (spc436_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 436, linebuf436);
          linebuf436 = "";
       end
    end else begin
       hitMadPrint436 = 0;
    end
  end
end


string linebuf437 = "";
logic hitMadPrint437 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc437_inst_done && ((spc437_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint437 = 1;
       linebuf437 = {linebuf437, spc437_phy_pc_w[8:1]};
       if (spc437_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 437, linebuf437);
          linebuf437 = "";
       end
    end else begin
       hitMadPrint437 = 0;
    end
  end
end


string linebuf438 = "";
logic hitMadPrint438 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc438_inst_done && ((spc438_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint438 = 1;
       linebuf438 = {linebuf438, spc438_phy_pc_w[8:1]};
       if (spc438_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 438, linebuf438);
          linebuf438 = "";
       end
    end else begin
       hitMadPrint438 = 0;
    end
  end
end


string linebuf439 = "";
logic hitMadPrint439 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc439_inst_done && ((spc439_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint439 = 1;
       linebuf439 = {linebuf439, spc439_phy_pc_w[8:1]};
       if (spc439_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 439, linebuf439);
          linebuf439 = "";
       end
    end else begin
       hitMadPrint439 = 0;
    end
  end
end


string linebuf440 = "";
logic hitMadPrint440 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc440_inst_done && ((spc440_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint440 = 1;
       linebuf440 = {linebuf440, spc440_phy_pc_w[8:1]};
       if (spc440_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 440, linebuf440);
          linebuf440 = "";
       end
    end else begin
       hitMadPrint440 = 0;
    end
  end
end


string linebuf441 = "";
logic hitMadPrint441 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc441_inst_done && ((spc441_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint441 = 1;
       linebuf441 = {linebuf441, spc441_phy_pc_w[8:1]};
       if (spc441_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 441, linebuf441);
          linebuf441 = "";
       end
    end else begin
       hitMadPrint441 = 0;
    end
  end
end


string linebuf442 = "";
logic hitMadPrint442 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc442_inst_done && ((spc442_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint442 = 1;
       linebuf442 = {linebuf442, spc442_phy_pc_w[8:1]};
       if (spc442_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 442, linebuf442);
          linebuf442 = "";
       end
    end else begin
       hitMadPrint442 = 0;
    end
  end
end


string linebuf443 = "";
logic hitMadPrint443 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc443_inst_done && ((spc443_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint443 = 1;
       linebuf443 = {linebuf443, spc443_phy_pc_w[8:1]};
       if (spc443_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 443, linebuf443);
          linebuf443 = "";
       end
    end else begin
       hitMadPrint443 = 0;
    end
  end
end


string linebuf444 = "";
logic hitMadPrint444 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc444_inst_done && ((spc444_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint444 = 1;
       linebuf444 = {linebuf444, spc444_phy_pc_w[8:1]};
       if (spc444_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 444, linebuf444);
          linebuf444 = "";
       end
    end else begin
       hitMadPrint444 = 0;
    end
  end
end


string linebuf445 = "";
logic hitMadPrint445 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc445_inst_done && ((spc445_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint445 = 1;
       linebuf445 = {linebuf445, spc445_phy_pc_w[8:1]};
       if (spc445_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 445, linebuf445);
          linebuf445 = "";
       end
    end else begin
       hitMadPrint445 = 0;
    end
  end
end


string linebuf446 = "";
logic hitMadPrint446 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc446_inst_done && ((spc446_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint446 = 1;
       linebuf446 = {linebuf446, spc446_phy_pc_w[8:1]};
       if (spc446_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 446, linebuf446);
          linebuf446 = "";
       end
    end else begin
       hitMadPrint446 = 0;
    end
  end
end


string linebuf447 = "";
logic hitMadPrint447 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc447_inst_done && ((spc447_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint447 = 1;
       linebuf447 = {linebuf447, spc447_phy_pc_w[8:1]};
       if (spc447_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 447, linebuf447);
          linebuf447 = "";
       end
    end else begin
       hitMadPrint447 = 0;
    end
  end
end


string linebuf448 = "";
logic hitMadPrint448 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc448_inst_done && ((spc448_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint448 = 1;
       linebuf448 = {linebuf448, spc448_phy_pc_w[8:1]};
       if (spc448_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 448, linebuf448);
          linebuf448 = "";
       end
    end else begin
       hitMadPrint448 = 0;
    end
  end
end


string linebuf449 = "";
logic hitMadPrint449 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc449_inst_done && ((spc449_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint449 = 1;
       linebuf449 = {linebuf449, spc449_phy_pc_w[8:1]};
       if (spc449_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 449, linebuf449);
          linebuf449 = "";
       end
    end else begin
       hitMadPrint449 = 0;
    end
  end
end


string linebuf450 = "";
logic hitMadPrint450 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc450_inst_done && ((spc450_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint450 = 1;
       linebuf450 = {linebuf450, spc450_phy_pc_w[8:1]};
       if (spc450_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 450, linebuf450);
          linebuf450 = "";
       end
    end else begin
       hitMadPrint450 = 0;
    end
  end
end


string linebuf451 = "";
logic hitMadPrint451 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc451_inst_done && ((spc451_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint451 = 1;
       linebuf451 = {linebuf451, spc451_phy_pc_w[8:1]};
       if (spc451_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 451, linebuf451);
          linebuf451 = "";
       end
    end else begin
       hitMadPrint451 = 0;
    end
  end
end


string linebuf452 = "";
logic hitMadPrint452 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc452_inst_done && ((spc452_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint452 = 1;
       linebuf452 = {linebuf452, spc452_phy_pc_w[8:1]};
       if (spc452_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 452, linebuf452);
          linebuf452 = "";
       end
    end else begin
       hitMadPrint452 = 0;
    end
  end
end


string linebuf453 = "";
logic hitMadPrint453 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc453_inst_done && ((spc453_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint453 = 1;
       linebuf453 = {linebuf453, spc453_phy_pc_w[8:1]};
       if (spc453_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 453, linebuf453);
          linebuf453 = "";
       end
    end else begin
       hitMadPrint453 = 0;
    end
  end
end


string linebuf454 = "";
logic hitMadPrint454 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc454_inst_done && ((spc454_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint454 = 1;
       linebuf454 = {linebuf454, spc454_phy_pc_w[8:1]};
       if (spc454_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 454, linebuf454);
          linebuf454 = "";
       end
    end else begin
       hitMadPrint454 = 0;
    end
  end
end


string linebuf455 = "";
logic hitMadPrint455 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc455_inst_done && ((spc455_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint455 = 1;
       linebuf455 = {linebuf455, spc455_phy_pc_w[8:1]};
       if (spc455_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 455, linebuf455);
          linebuf455 = "";
       end
    end else begin
       hitMadPrint455 = 0;
    end
  end
end


string linebuf456 = "";
logic hitMadPrint456 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc456_inst_done && ((spc456_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint456 = 1;
       linebuf456 = {linebuf456, spc456_phy_pc_w[8:1]};
       if (spc456_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 456, linebuf456);
          linebuf456 = "";
       end
    end else begin
       hitMadPrint456 = 0;
    end
  end
end


string linebuf457 = "";
logic hitMadPrint457 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc457_inst_done && ((spc457_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint457 = 1;
       linebuf457 = {linebuf457, spc457_phy_pc_w[8:1]};
       if (spc457_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 457, linebuf457);
          linebuf457 = "";
       end
    end else begin
       hitMadPrint457 = 0;
    end
  end
end


string linebuf458 = "";
logic hitMadPrint458 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc458_inst_done && ((spc458_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint458 = 1;
       linebuf458 = {linebuf458, spc458_phy_pc_w[8:1]};
       if (spc458_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 458, linebuf458);
          linebuf458 = "";
       end
    end else begin
       hitMadPrint458 = 0;
    end
  end
end


string linebuf459 = "";
logic hitMadPrint459 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc459_inst_done && ((spc459_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint459 = 1;
       linebuf459 = {linebuf459, spc459_phy_pc_w[8:1]};
       if (spc459_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 459, linebuf459);
          linebuf459 = "";
       end
    end else begin
       hitMadPrint459 = 0;
    end
  end
end


string linebuf460 = "";
logic hitMadPrint460 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc460_inst_done && ((spc460_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint460 = 1;
       linebuf460 = {linebuf460, spc460_phy_pc_w[8:1]};
       if (spc460_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 460, linebuf460);
          linebuf460 = "";
       end
    end else begin
       hitMadPrint460 = 0;
    end
  end
end


string linebuf461 = "";
logic hitMadPrint461 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc461_inst_done && ((spc461_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint461 = 1;
       linebuf461 = {linebuf461, spc461_phy_pc_w[8:1]};
       if (spc461_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 461, linebuf461);
          linebuf461 = "";
       end
    end else begin
       hitMadPrint461 = 0;
    end
  end
end


string linebuf462 = "";
logic hitMadPrint462 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc462_inst_done && ((spc462_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint462 = 1;
       linebuf462 = {linebuf462, spc462_phy_pc_w[8:1]};
       if (spc462_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 462, linebuf462);
          linebuf462 = "";
       end
    end else begin
       hitMadPrint462 = 0;
    end
  end
end


string linebuf463 = "";
logic hitMadPrint463 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc463_inst_done && ((spc463_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint463 = 1;
       linebuf463 = {linebuf463, spc463_phy_pc_w[8:1]};
       if (spc463_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 463, linebuf463);
          linebuf463 = "";
       end
    end else begin
       hitMadPrint463 = 0;
    end
  end
end


string linebuf464 = "";
logic hitMadPrint464 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc464_inst_done && ((spc464_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint464 = 1;
       linebuf464 = {linebuf464, spc464_phy_pc_w[8:1]};
       if (spc464_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 464, linebuf464);
          linebuf464 = "";
       end
    end else begin
       hitMadPrint464 = 0;
    end
  end
end


string linebuf465 = "";
logic hitMadPrint465 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc465_inst_done && ((spc465_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint465 = 1;
       linebuf465 = {linebuf465, spc465_phy_pc_w[8:1]};
       if (spc465_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 465, linebuf465);
          linebuf465 = "";
       end
    end else begin
       hitMadPrint465 = 0;
    end
  end
end


string linebuf466 = "";
logic hitMadPrint466 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc466_inst_done && ((spc466_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint466 = 1;
       linebuf466 = {linebuf466, spc466_phy_pc_w[8:1]};
       if (spc466_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 466, linebuf466);
          linebuf466 = "";
       end
    end else begin
       hitMadPrint466 = 0;
    end
  end
end


string linebuf467 = "";
logic hitMadPrint467 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc467_inst_done && ((spc467_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint467 = 1;
       linebuf467 = {linebuf467, spc467_phy_pc_w[8:1]};
       if (spc467_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 467, linebuf467);
          linebuf467 = "";
       end
    end else begin
       hitMadPrint467 = 0;
    end
  end
end


string linebuf468 = "";
logic hitMadPrint468 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc468_inst_done && ((spc468_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint468 = 1;
       linebuf468 = {linebuf468, spc468_phy_pc_w[8:1]};
       if (spc468_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 468, linebuf468);
          linebuf468 = "";
       end
    end else begin
       hitMadPrint468 = 0;
    end
  end
end


string linebuf469 = "";
logic hitMadPrint469 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc469_inst_done && ((spc469_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint469 = 1;
       linebuf469 = {linebuf469, spc469_phy_pc_w[8:1]};
       if (spc469_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 469, linebuf469);
          linebuf469 = "";
       end
    end else begin
       hitMadPrint469 = 0;
    end
  end
end


string linebuf470 = "";
logic hitMadPrint470 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc470_inst_done && ((spc470_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint470 = 1;
       linebuf470 = {linebuf470, spc470_phy_pc_w[8:1]};
       if (spc470_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 470, linebuf470);
          linebuf470 = "";
       end
    end else begin
       hitMadPrint470 = 0;
    end
  end
end


string linebuf471 = "";
logic hitMadPrint471 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc471_inst_done && ((spc471_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint471 = 1;
       linebuf471 = {linebuf471, spc471_phy_pc_w[8:1]};
       if (spc471_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 471, linebuf471);
          linebuf471 = "";
       end
    end else begin
       hitMadPrint471 = 0;
    end
  end
end


string linebuf472 = "";
logic hitMadPrint472 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc472_inst_done && ((spc472_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint472 = 1;
       linebuf472 = {linebuf472, spc472_phy_pc_w[8:1]};
       if (spc472_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 472, linebuf472);
          linebuf472 = "";
       end
    end else begin
       hitMadPrint472 = 0;
    end
  end
end


string linebuf473 = "";
logic hitMadPrint473 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc473_inst_done && ((spc473_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint473 = 1;
       linebuf473 = {linebuf473, spc473_phy_pc_w[8:1]};
       if (spc473_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 473, linebuf473);
          linebuf473 = "";
       end
    end else begin
       hitMadPrint473 = 0;
    end
  end
end


string linebuf474 = "";
logic hitMadPrint474 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc474_inst_done && ((spc474_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint474 = 1;
       linebuf474 = {linebuf474, spc474_phy_pc_w[8:1]};
       if (spc474_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 474, linebuf474);
          linebuf474 = "";
       end
    end else begin
       hitMadPrint474 = 0;
    end
  end
end


string linebuf475 = "";
logic hitMadPrint475 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc475_inst_done && ((spc475_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint475 = 1;
       linebuf475 = {linebuf475, spc475_phy_pc_w[8:1]};
       if (spc475_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 475, linebuf475);
          linebuf475 = "";
       end
    end else begin
       hitMadPrint475 = 0;
    end
  end
end


string linebuf476 = "";
logic hitMadPrint476 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc476_inst_done && ((spc476_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint476 = 1;
       linebuf476 = {linebuf476, spc476_phy_pc_w[8:1]};
       if (spc476_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 476, linebuf476);
          linebuf476 = "";
       end
    end else begin
       hitMadPrint476 = 0;
    end
  end
end


string linebuf477 = "";
logic hitMadPrint477 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc477_inst_done && ((spc477_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint477 = 1;
       linebuf477 = {linebuf477, spc477_phy_pc_w[8:1]};
       if (spc477_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 477, linebuf477);
          linebuf477 = "";
       end
    end else begin
       hitMadPrint477 = 0;
    end
  end
end


string linebuf478 = "";
logic hitMadPrint478 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc478_inst_done && ((spc478_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint478 = 1;
       linebuf478 = {linebuf478, spc478_phy_pc_w[8:1]};
       if (spc478_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 478, linebuf478);
          linebuf478 = "";
       end
    end else begin
       hitMadPrint478 = 0;
    end
  end
end


string linebuf479 = "";
logic hitMadPrint479 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc479_inst_done && ((spc479_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint479 = 1;
       linebuf479 = {linebuf479, spc479_phy_pc_w[8:1]};
       if (spc479_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 479, linebuf479);
          linebuf479 = "";
       end
    end else begin
       hitMadPrint479 = 0;
    end
  end
end


string linebuf480 = "";
logic hitMadPrint480 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc480_inst_done && ((spc480_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint480 = 1;
       linebuf480 = {linebuf480, spc480_phy_pc_w[8:1]};
       if (spc480_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 480, linebuf480);
          linebuf480 = "";
       end
    end else begin
       hitMadPrint480 = 0;
    end
  end
end


string linebuf481 = "";
logic hitMadPrint481 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc481_inst_done && ((spc481_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint481 = 1;
       linebuf481 = {linebuf481, spc481_phy_pc_w[8:1]};
       if (spc481_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 481, linebuf481);
          linebuf481 = "";
       end
    end else begin
       hitMadPrint481 = 0;
    end
  end
end


string linebuf482 = "";
logic hitMadPrint482 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc482_inst_done && ((spc482_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint482 = 1;
       linebuf482 = {linebuf482, spc482_phy_pc_w[8:1]};
       if (spc482_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 482, linebuf482);
          linebuf482 = "";
       end
    end else begin
       hitMadPrint482 = 0;
    end
  end
end


string linebuf483 = "";
logic hitMadPrint483 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc483_inst_done && ((spc483_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint483 = 1;
       linebuf483 = {linebuf483, spc483_phy_pc_w[8:1]};
       if (spc483_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 483, linebuf483);
          linebuf483 = "";
       end
    end else begin
       hitMadPrint483 = 0;
    end
  end
end


string linebuf484 = "";
logic hitMadPrint484 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc484_inst_done && ((spc484_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint484 = 1;
       linebuf484 = {linebuf484, spc484_phy_pc_w[8:1]};
       if (spc484_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 484, linebuf484);
          linebuf484 = "";
       end
    end else begin
       hitMadPrint484 = 0;
    end
  end
end


string linebuf485 = "";
logic hitMadPrint485 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc485_inst_done && ((spc485_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint485 = 1;
       linebuf485 = {linebuf485, spc485_phy_pc_w[8:1]};
       if (spc485_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 485, linebuf485);
          linebuf485 = "";
       end
    end else begin
       hitMadPrint485 = 0;
    end
  end
end


string linebuf486 = "";
logic hitMadPrint486 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc486_inst_done && ((spc486_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint486 = 1;
       linebuf486 = {linebuf486, spc486_phy_pc_w[8:1]};
       if (spc486_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 486, linebuf486);
          linebuf486 = "";
       end
    end else begin
       hitMadPrint486 = 0;
    end
  end
end


string linebuf487 = "";
logic hitMadPrint487 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc487_inst_done && ((spc487_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint487 = 1;
       linebuf487 = {linebuf487, spc487_phy_pc_w[8:1]};
       if (spc487_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 487, linebuf487);
          linebuf487 = "";
       end
    end else begin
       hitMadPrint487 = 0;
    end
  end
end


string linebuf488 = "";
logic hitMadPrint488 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc488_inst_done && ((spc488_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint488 = 1;
       linebuf488 = {linebuf488, spc488_phy_pc_w[8:1]};
       if (spc488_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 488, linebuf488);
          linebuf488 = "";
       end
    end else begin
       hitMadPrint488 = 0;
    end
  end
end


string linebuf489 = "";
logic hitMadPrint489 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc489_inst_done && ((spc489_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint489 = 1;
       linebuf489 = {linebuf489, spc489_phy_pc_w[8:1]};
       if (spc489_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 489, linebuf489);
          linebuf489 = "";
       end
    end else begin
       hitMadPrint489 = 0;
    end
  end
end


string linebuf490 = "";
logic hitMadPrint490 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc490_inst_done && ((spc490_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint490 = 1;
       linebuf490 = {linebuf490, spc490_phy_pc_w[8:1]};
       if (spc490_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 490, linebuf490);
          linebuf490 = "";
       end
    end else begin
       hitMadPrint490 = 0;
    end
  end
end


string linebuf491 = "";
logic hitMadPrint491 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc491_inst_done && ((spc491_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint491 = 1;
       linebuf491 = {linebuf491, spc491_phy_pc_w[8:1]};
       if (spc491_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 491, linebuf491);
          linebuf491 = "";
       end
    end else begin
       hitMadPrint491 = 0;
    end
  end
end


string linebuf492 = "";
logic hitMadPrint492 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc492_inst_done && ((spc492_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint492 = 1;
       linebuf492 = {linebuf492, spc492_phy_pc_w[8:1]};
       if (spc492_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 492, linebuf492);
          linebuf492 = "";
       end
    end else begin
       hitMadPrint492 = 0;
    end
  end
end


string linebuf493 = "";
logic hitMadPrint493 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc493_inst_done && ((spc493_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint493 = 1;
       linebuf493 = {linebuf493, spc493_phy_pc_w[8:1]};
       if (spc493_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 493, linebuf493);
          linebuf493 = "";
       end
    end else begin
       hitMadPrint493 = 0;
    end
  end
end


string linebuf494 = "";
logic hitMadPrint494 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc494_inst_done && ((spc494_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint494 = 1;
       linebuf494 = {linebuf494, spc494_phy_pc_w[8:1]};
       if (spc494_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 494, linebuf494);
          linebuf494 = "";
       end
    end else begin
       hitMadPrint494 = 0;
    end
  end
end


string linebuf495 = "";
logic hitMadPrint495 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc495_inst_done && ((spc495_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint495 = 1;
       linebuf495 = {linebuf495, spc495_phy_pc_w[8:1]};
       if (spc495_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 495, linebuf495);
          linebuf495 = "";
       end
    end else begin
       hitMadPrint495 = 0;
    end
  end
end


string linebuf496 = "";
logic hitMadPrint496 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc496_inst_done && ((spc496_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint496 = 1;
       linebuf496 = {linebuf496, spc496_phy_pc_w[8:1]};
       if (spc496_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 496, linebuf496);
          linebuf496 = "";
       end
    end else begin
       hitMadPrint496 = 0;
    end
  end
end


string linebuf497 = "";
logic hitMadPrint497 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc497_inst_done && ((spc497_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint497 = 1;
       linebuf497 = {linebuf497, spc497_phy_pc_w[8:1]};
       if (spc497_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 497, linebuf497);
          linebuf497 = "";
       end
    end else begin
       hitMadPrint497 = 0;
    end
  end
end


string linebuf498 = "";
logic hitMadPrint498 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc498_inst_done && ((spc498_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint498 = 1;
       linebuf498 = {linebuf498, spc498_phy_pc_w[8:1]};
       if (spc498_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 498, linebuf498);
          linebuf498 = "";
       end
    end else begin
       hitMadPrint498 = 0;
    end
  end
end


string linebuf499 = "";
logic hitMadPrint499 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc499_inst_done && ((spc499_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint499 = 1;
       linebuf499 = {linebuf499, spc499_phy_pc_w[8:1]};
       if (spc499_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 499, linebuf499);
          linebuf499 = "";
       end
    end else begin
       hitMadPrint499 = 0;
    end
  end
end


string linebuf500 = "";
logic hitMadPrint500 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc500_inst_done && ((spc500_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint500 = 1;
       linebuf500 = {linebuf500, spc500_phy_pc_w[8:1]};
       if (spc500_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 500, linebuf500);
          linebuf500 = "";
       end
    end else begin
       hitMadPrint500 = 0;
    end
  end
end


string linebuf501 = "";
logic hitMadPrint501 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc501_inst_done && ((spc501_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint501 = 1;
       linebuf501 = {linebuf501, spc501_phy_pc_w[8:1]};
       if (spc501_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 501, linebuf501);
          linebuf501 = "";
       end
    end else begin
       hitMadPrint501 = 0;
    end
  end
end


string linebuf502 = "";
logic hitMadPrint502 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc502_inst_done && ((spc502_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint502 = 1;
       linebuf502 = {linebuf502, spc502_phy_pc_w[8:1]};
       if (spc502_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 502, linebuf502);
          linebuf502 = "";
       end
    end else begin
       hitMadPrint502 = 0;
    end
  end
end


string linebuf503 = "";
logic hitMadPrint503 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc503_inst_done && ((spc503_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint503 = 1;
       linebuf503 = {linebuf503, spc503_phy_pc_w[8:1]};
       if (spc503_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 503, linebuf503);
          linebuf503 = "";
       end
    end else begin
       hitMadPrint503 = 0;
    end
  end
end


string linebuf504 = "";
logic hitMadPrint504 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc504_inst_done && ((spc504_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint504 = 1;
       linebuf504 = {linebuf504, spc504_phy_pc_w[8:1]};
       if (spc504_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 504, linebuf504);
          linebuf504 = "";
       end
    end else begin
       hitMadPrint504 = 0;
    end
  end
end


string linebuf505 = "";
logic hitMadPrint505 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc505_inst_done && ((spc505_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint505 = 1;
       linebuf505 = {linebuf505, spc505_phy_pc_w[8:1]};
       if (spc505_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 505, linebuf505);
          linebuf505 = "";
       end
    end else begin
       hitMadPrint505 = 0;
    end
  end
end


string linebuf506 = "";
logic hitMadPrint506 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc506_inst_done && ((spc506_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint506 = 1;
       linebuf506 = {linebuf506, spc506_phy_pc_w[8:1]};
       if (spc506_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 506, linebuf506);
          linebuf506 = "";
       end
    end else begin
       hitMadPrint506 = 0;
    end
  end
end


string linebuf507 = "";
logic hitMadPrint507 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc507_inst_done && ((spc507_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint507 = 1;
       linebuf507 = {linebuf507, spc507_phy_pc_w[8:1]};
       if (spc507_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 507, linebuf507);
          linebuf507 = "";
       end
    end else begin
       hitMadPrint507 = 0;
    end
  end
end


string linebuf508 = "";
logic hitMadPrint508 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc508_inst_done && ((spc508_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint508 = 1;
       linebuf508 = {linebuf508, spc508_phy_pc_w[8:1]};
       if (spc508_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 508, linebuf508);
          linebuf508 = "";
       end
    end else begin
       hitMadPrint508 = 0;
    end
  end
end


string linebuf509 = "";
logic hitMadPrint509 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc509_inst_done && ((spc509_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint509 = 1;
       linebuf509 = {linebuf509, spc509_phy_pc_w[8:1]};
       if (spc509_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 509, linebuf509);
          linebuf509 = "";
       end
    end else begin
       hitMadPrint509 = 0;
    end
  end
end


string linebuf510 = "";
logic hitMadPrint510 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc510_inst_done && ((spc510_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint510 = 1;
       linebuf510 = {linebuf510, spc510_phy_pc_w[8:1]};
       if (spc510_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 510, linebuf510);
          linebuf510 = "";
       end
    end else begin
       hitMadPrint510 = 0;
    end
  end
end


string linebuf511 = "";
logic hitMadPrint511 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc511_inst_done && ((spc511_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint511 = 1;
       linebuf511 = {linebuf511, spc511_phy_pc_w[8:1]};
       if (spc511_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 511, linebuf511);
          linebuf511 = "";
       end
    end else begin
       hitMadPrint511 = 0;
    end
  end
end


string linebuf512 = "";
logic hitMadPrint512 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc512_inst_done && ((spc512_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint512 = 1;
       linebuf512 = {linebuf512, spc512_phy_pc_w[8:1]};
       if (spc512_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 512, linebuf512);
          linebuf512 = "";
       end
    end else begin
       hitMadPrint512 = 0;
    end
  end
end


string linebuf513 = "";
logic hitMadPrint513 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc513_inst_done && ((spc513_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint513 = 1;
       linebuf513 = {linebuf513, spc513_phy_pc_w[8:1]};
       if (spc513_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 513, linebuf513);
          linebuf513 = "";
       end
    end else begin
       hitMadPrint513 = 0;
    end
  end
end


string linebuf514 = "";
logic hitMadPrint514 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc514_inst_done && ((spc514_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint514 = 1;
       linebuf514 = {linebuf514, spc514_phy_pc_w[8:1]};
       if (spc514_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 514, linebuf514);
          linebuf514 = "";
       end
    end else begin
       hitMadPrint514 = 0;
    end
  end
end


string linebuf515 = "";
logic hitMadPrint515 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc515_inst_done && ((spc515_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint515 = 1;
       linebuf515 = {linebuf515, spc515_phy_pc_w[8:1]};
       if (spc515_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 515, linebuf515);
          linebuf515 = "";
       end
    end else begin
       hitMadPrint515 = 0;
    end
  end
end


string linebuf516 = "";
logic hitMadPrint516 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc516_inst_done && ((spc516_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint516 = 1;
       linebuf516 = {linebuf516, spc516_phy_pc_w[8:1]};
       if (spc516_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 516, linebuf516);
          linebuf516 = "";
       end
    end else begin
       hitMadPrint516 = 0;
    end
  end
end


string linebuf517 = "";
logic hitMadPrint517 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc517_inst_done && ((spc517_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint517 = 1;
       linebuf517 = {linebuf517, spc517_phy_pc_w[8:1]};
       if (spc517_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 517, linebuf517);
          linebuf517 = "";
       end
    end else begin
       hitMadPrint517 = 0;
    end
  end
end


string linebuf518 = "";
logic hitMadPrint518 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc518_inst_done && ((spc518_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint518 = 1;
       linebuf518 = {linebuf518, spc518_phy_pc_w[8:1]};
       if (spc518_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 518, linebuf518);
          linebuf518 = "";
       end
    end else begin
       hitMadPrint518 = 0;
    end
  end
end


string linebuf519 = "";
logic hitMadPrint519 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc519_inst_done && ((spc519_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint519 = 1;
       linebuf519 = {linebuf519, spc519_phy_pc_w[8:1]};
       if (spc519_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 519, linebuf519);
          linebuf519 = "";
       end
    end else begin
       hitMadPrint519 = 0;
    end
  end
end


string linebuf520 = "";
logic hitMadPrint520 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc520_inst_done && ((spc520_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint520 = 1;
       linebuf520 = {linebuf520, spc520_phy_pc_w[8:1]};
       if (spc520_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 520, linebuf520);
          linebuf520 = "";
       end
    end else begin
       hitMadPrint520 = 0;
    end
  end
end


string linebuf521 = "";
logic hitMadPrint521 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc521_inst_done && ((spc521_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint521 = 1;
       linebuf521 = {linebuf521, spc521_phy_pc_w[8:1]};
       if (spc521_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 521, linebuf521);
          linebuf521 = "";
       end
    end else begin
       hitMadPrint521 = 0;
    end
  end
end


string linebuf522 = "";
logic hitMadPrint522 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc522_inst_done && ((spc522_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint522 = 1;
       linebuf522 = {linebuf522, spc522_phy_pc_w[8:1]};
       if (spc522_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 522, linebuf522);
          linebuf522 = "";
       end
    end else begin
       hitMadPrint522 = 0;
    end
  end
end


string linebuf523 = "";
logic hitMadPrint523 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc523_inst_done && ((spc523_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint523 = 1;
       linebuf523 = {linebuf523, spc523_phy_pc_w[8:1]};
       if (spc523_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 523, linebuf523);
          linebuf523 = "";
       end
    end else begin
       hitMadPrint523 = 0;
    end
  end
end


string linebuf524 = "";
logic hitMadPrint524 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc524_inst_done && ((spc524_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint524 = 1;
       linebuf524 = {linebuf524, spc524_phy_pc_w[8:1]};
       if (spc524_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 524, linebuf524);
          linebuf524 = "";
       end
    end else begin
       hitMadPrint524 = 0;
    end
  end
end


string linebuf525 = "";
logic hitMadPrint525 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc525_inst_done && ((spc525_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint525 = 1;
       linebuf525 = {linebuf525, spc525_phy_pc_w[8:1]};
       if (spc525_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 525, linebuf525);
          linebuf525 = "";
       end
    end else begin
       hitMadPrint525 = 0;
    end
  end
end


string linebuf526 = "";
logic hitMadPrint526 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc526_inst_done && ((spc526_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint526 = 1;
       linebuf526 = {linebuf526, spc526_phy_pc_w[8:1]};
       if (spc526_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 526, linebuf526);
          linebuf526 = "";
       end
    end else begin
       hitMadPrint526 = 0;
    end
  end
end


string linebuf527 = "";
logic hitMadPrint527 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc527_inst_done && ((spc527_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint527 = 1;
       linebuf527 = {linebuf527, spc527_phy_pc_w[8:1]};
       if (spc527_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 527, linebuf527);
          linebuf527 = "";
       end
    end else begin
       hitMadPrint527 = 0;
    end
  end
end


string linebuf528 = "";
logic hitMadPrint528 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc528_inst_done && ((spc528_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint528 = 1;
       linebuf528 = {linebuf528, spc528_phy_pc_w[8:1]};
       if (spc528_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 528, linebuf528);
          linebuf528 = "";
       end
    end else begin
       hitMadPrint528 = 0;
    end
  end
end


string linebuf529 = "";
logic hitMadPrint529 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc529_inst_done && ((spc529_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint529 = 1;
       linebuf529 = {linebuf529, spc529_phy_pc_w[8:1]};
       if (spc529_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 529, linebuf529);
          linebuf529 = "";
       end
    end else begin
       hitMadPrint529 = 0;
    end
  end
end


string linebuf530 = "";
logic hitMadPrint530 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc530_inst_done && ((spc530_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint530 = 1;
       linebuf530 = {linebuf530, spc530_phy_pc_w[8:1]};
       if (spc530_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 530, linebuf530);
          linebuf530 = "";
       end
    end else begin
       hitMadPrint530 = 0;
    end
  end
end


string linebuf531 = "";
logic hitMadPrint531 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc531_inst_done && ((spc531_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint531 = 1;
       linebuf531 = {linebuf531, spc531_phy_pc_w[8:1]};
       if (spc531_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 531, linebuf531);
          linebuf531 = "";
       end
    end else begin
       hitMadPrint531 = 0;
    end
  end
end


string linebuf532 = "";
logic hitMadPrint532 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc532_inst_done && ((spc532_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint532 = 1;
       linebuf532 = {linebuf532, spc532_phy_pc_w[8:1]};
       if (spc532_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 532, linebuf532);
          linebuf532 = "";
       end
    end else begin
       hitMadPrint532 = 0;
    end
  end
end


string linebuf533 = "";
logic hitMadPrint533 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc533_inst_done && ((spc533_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint533 = 1;
       linebuf533 = {linebuf533, spc533_phy_pc_w[8:1]};
       if (spc533_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 533, linebuf533);
          linebuf533 = "";
       end
    end else begin
       hitMadPrint533 = 0;
    end
  end
end


string linebuf534 = "";
logic hitMadPrint534 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc534_inst_done && ((spc534_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint534 = 1;
       linebuf534 = {linebuf534, spc534_phy_pc_w[8:1]};
       if (spc534_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 534, linebuf534);
          linebuf534 = "";
       end
    end else begin
       hitMadPrint534 = 0;
    end
  end
end


string linebuf535 = "";
logic hitMadPrint535 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc535_inst_done && ((spc535_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint535 = 1;
       linebuf535 = {linebuf535, spc535_phy_pc_w[8:1]};
       if (spc535_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 535, linebuf535);
          linebuf535 = "";
       end
    end else begin
       hitMadPrint535 = 0;
    end
  end
end


string linebuf536 = "";
logic hitMadPrint536 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc536_inst_done && ((spc536_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint536 = 1;
       linebuf536 = {linebuf536, spc536_phy_pc_w[8:1]};
       if (spc536_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 536, linebuf536);
          linebuf536 = "";
       end
    end else begin
       hitMadPrint536 = 0;
    end
  end
end


string linebuf537 = "";
logic hitMadPrint537 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc537_inst_done && ((spc537_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint537 = 1;
       linebuf537 = {linebuf537, spc537_phy_pc_w[8:1]};
       if (spc537_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 537, linebuf537);
          linebuf537 = "";
       end
    end else begin
       hitMadPrint537 = 0;
    end
  end
end


string linebuf538 = "";
logic hitMadPrint538 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc538_inst_done && ((spc538_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint538 = 1;
       linebuf538 = {linebuf538, spc538_phy_pc_w[8:1]};
       if (spc538_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 538, linebuf538);
          linebuf538 = "";
       end
    end else begin
       hitMadPrint538 = 0;
    end
  end
end


string linebuf539 = "";
logic hitMadPrint539 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc539_inst_done && ((spc539_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint539 = 1;
       linebuf539 = {linebuf539, spc539_phy_pc_w[8:1]};
       if (spc539_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 539, linebuf539);
          linebuf539 = "";
       end
    end else begin
       hitMadPrint539 = 0;
    end
  end
end


string linebuf540 = "";
logic hitMadPrint540 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc540_inst_done && ((spc540_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint540 = 1;
       linebuf540 = {linebuf540, spc540_phy_pc_w[8:1]};
       if (spc540_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 540, linebuf540);
          linebuf540 = "";
       end
    end else begin
       hitMadPrint540 = 0;
    end
  end
end


string linebuf541 = "";
logic hitMadPrint541 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc541_inst_done && ((spc541_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint541 = 1;
       linebuf541 = {linebuf541, spc541_phy_pc_w[8:1]};
       if (spc541_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 541, linebuf541);
          linebuf541 = "";
       end
    end else begin
       hitMadPrint541 = 0;
    end
  end
end


string linebuf542 = "";
logic hitMadPrint542 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc542_inst_done && ((spc542_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint542 = 1;
       linebuf542 = {linebuf542, spc542_phy_pc_w[8:1]};
       if (spc542_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 542, linebuf542);
          linebuf542 = "";
       end
    end else begin
       hitMadPrint542 = 0;
    end
  end
end


string linebuf543 = "";
logic hitMadPrint543 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc543_inst_done && ((spc543_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint543 = 1;
       linebuf543 = {linebuf543, spc543_phy_pc_w[8:1]};
       if (spc543_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 543, linebuf543);
          linebuf543 = "";
       end
    end else begin
       hitMadPrint543 = 0;
    end
  end
end


string linebuf544 = "";
logic hitMadPrint544 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc544_inst_done && ((spc544_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint544 = 1;
       linebuf544 = {linebuf544, spc544_phy_pc_w[8:1]};
       if (spc544_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 544, linebuf544);
          linebuf544 = "";
       end
    end else begin
       hitMadPrint544 = 0;
    end
  end
end


string linebuf545 = "";
logic hitMadPrint545 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc545_inst_done && ((spc545_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint545 = 1;
       linebuf545 = {linebuf545, spc545_phy_pc_w[8:1]};
       if (spc545_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 545, linebuf545);
          linebuf545 = "";
       end
    end else begin
       hitMadPrint545 = 0;
    end
  end
end


string linebuf546 = "";
logic hitMadPrint546 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc546_inst_done && ((spc546_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint546 = 1;
       linebuf546 = {linebuf546, spc546_phy_pc_w[8:1]};
       if (spc546_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 546, linebuf546);
          linebuf546 = "";
       end
    end else begin
       hitMadPrint546 = 0;
    end
  end
end


string linebuf547 = "";
logic hitMadPrint547 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc547_inst_done && ((spc547_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint547 = 1;
       linebuf547 = {linebuf547, spc547_phy_pc_w[8:1]};
       if (spc547_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 547, linebuf547);
          linebuf547 = "";
       end
    end else begin
       hitMadPrint547 = 0;
    end
  end
end


string linebuf548 = "";
logic hitMadPrint548 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc548_inst_done && ((spc548_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint548 = 1;
       linebuf548 = {linebuf548, spc548_phy_pc_w[8:1]};
       if (spc548_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 548, linebuf548);
          linebuf548 = "";
       end
    end else begin
       hitMadPrint548 = 0;
    end
  end
end


string linebuf549 = "";
logic hitMadPrint549 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc549_inst_done && ((spc549_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint549 = 1;
       linebuf549 = {linebuf549, spc549_phy_pc_w[8:1]};
       if (spc549_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 549, linebuf549);
          linebuf549 = "";
       end
    end else begin
       hitMadPrint549 = 0;
    end
  end
end


string linebuf550 = "";
logic hitMadPrint550 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc550_inst_done && ((spc550_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint550 = 1;
       linebuf550 = {linebuf550, spc550_phy_pc_w[8:1]};
       if (spc550_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 550, linebuf550);
          linebuf550 = "";
       end
    end else begin
       hitMadPrint550 = 0;
    end
  end
end


string linebuf551 = "";
logic hitMadPrint551 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc551_inst_done && ((spc551_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint551 = 1;
       linebuf551 = {linebuf551, spc551_phy_pc_w[8:1]};
       if (spc551_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 551, linebuf551);
          linebuf551 = "";
       end
    end else begin
       hitMadPrint551 = 0;
    end
  end
end


string linebuf552 = "";
logic hitMadPrint552 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc552_inst_done && ((spc552_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint552 = 1;
       linebuf552 = {linebuf552, spc552_phy_pc_w[8:1]};
       if (spc552_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 552, linebuf552);
          linebuf552 = "";
       end
    end else begin
       hitMadPrint552 = 0;
    end
  end
end


string linebuf553 = "";
logic hitMadPrint553 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc553_inst_done && ((spc553_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint553 = 1;
       linebuf553 = {linebuf553, spc553_phy_pc_w[8:1]};
       if (spc553_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 553, linebuf553);
          linebuf553 = "";
       end
    end else begin
       hitMadPrint553 = 0;
    end
  end
end


string linebuf554 = "";
logic hitMadPrint554 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc554_inst_done && ((spc554_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint554 = 1;
       linebuf554 = {linebuf554, spc554_phy_pc_w[8:1]};
       if (spc554_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 554, linebuf554);
          linebuf554 = "";
       end
    end else begin
       hitMadPrint554 = 0;
    end
  end
end


string linebuf555 = "";
logic hitMadPrint555 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc555_inst_done && ((spc555_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint555 = 1;
       linebuf555 = {linebuf555, spc555_phy_pc_w[8:1]};
       if (spc555_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 555, linebuf555);
          linebuf555 = "";
       end
    end else begin
       hitMadPrint555 = 0;
    end
  end
end


string linebuf556 = "";
logic hitMadPrint556 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc556_inst_done && ((spc556_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint556 = 1;
       linebuf556 = {linebuf556, spc556_phy_pc_w[8:1]};
       if (spc556_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 556, linebuf556);
          linebuf556 = "";
       end
    end else begin
       hitMadPrint556 = 0;
    end
  end
end


string linebuf557 = "";
logic hitMadPrint557 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc557_inst_done && ((spc557_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint557 = 1;
       linebuf557 = {linebuf557, spc557_phy_pc_w[8:1]};
       if (spc557_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 557, linebuf557);
          linebuf557 = "";
       end
    end else begin
       hitMadPrint557 = 0;
    end
  end
end


string linebuf558 = "";
logic hitMadPrint558 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc558_inst_done && ((spc558_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint558 = 1;
       linebuf558 = {linebuf558, spc558_phy_pc_w[8:1]};
       if (spc558_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 558, linebuf558);
          linebuf558 = "";
       end
    end else begin
       hitMadPrint558 = 0;
    end
  end
end


string linebuf559 = "";
logic hitMadPrint559 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc559_inst_done && ((spc559_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint559 = 1;
       linebuf559 = {linebuf559, spc559_phy_pc_w[8:1]};
       if (spc559_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 559, linebuf559);
          linebuf559 = "";
       end
    end else begin
       hitMadPrint559 = 0;
    end
  end
end


string linebuf560 = "";
logic hitMadPrint560 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc560_inst_done && ((spc560_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint560 = 1;
       linebuf560 = {linebuf560, spc560_phy_pc_w[8:1]};
       if (spc560_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 560, linebuf560);
          linebuf560 = "";
       end
    end else begin
       hitMadPrint560 = 0;
    end
  end
end


string linebuf561 = "";
logic hitMadPrint561 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc561_inst_done && ((spc561_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint561 = 1;
       linebuf561 = {linebuf561, spc561_phy_pc_w[8:1]};
       if (spc561_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 561, linebuf561);
          linebuf561 = "";
       end
    end else begin
       hitMadPrint561 = 0;
    end
  end
end


string linebuf562 = "";
logic hitMadPrint562 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc562_inst_done && ((spc562_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint562 = 1;
       linebuf562 = {linebuf562, spc562_phy_pc_w[8:1]};
       if (spc562_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 562, linebuf562);
          linebuf562 = "";
       end
    end else begin
       hitMadPrint562 = 0;
    end
  end
end


string linebuf563 = "";
logic hitMadPrint563 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc563_inst_done && ((spc563_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint563 = 1;
       linebuf563 = {linebuf563, spc563_phy_pc_w[8:1]};
       if (spc563_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 563, linebuf563);
          linebuf563 = "";
       end
    end else begin
       hitMadPrint563 = 0;
    end
  end
end


string linebuf564 = "";
logic hitMadPrint564 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc564_inst_done && ((spc564_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint564 = 1;
       linebuf564 = {linebuf564, spc564_phy_pc_w[8:1]};
       if (spc564_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 564, linebuf564);
          linebuf564 = "";
       end
    end else begin
       hitMadPrint564 = 0;
    end
  end
end


string linebuf565 = "";
logic hitMadPrint565 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc565_inst_done && ((spc565_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint565 = 1;
       linebuf565 = {linebuf565, spc565_phy_pc_w[8:1]};
       if (spc565_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 565, linebuf565);
          linebuf565 = "";
       end
    end else begin
       hitMadPrint565 = 0;
    end
  end
end


string linebuf566 = "";
logic hitMadPrint566 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc566_inst_done && ((spc566_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint566 = 1;
       linebuf566 = {linebuf566, spc566_phy_pc_w[8:1]};
       if (spc566_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 566, linebuf566);
          linebuf566 = "";
       end
    end else begin
       hitMadPrint566 = 0;
    end
  end
end


string linebuf567 = "";
logic hitMadPrint567 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc567_inst_done && ((spc567_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint567 = 1;
       linebuf567 = {linebuf567, spc567_phy_pc_w[8:1]};
       if (spc567_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 567, linebuf567);
          linebuf567 = "";
       end
    end else begin
       hitMadPrint567 = 0;
    end
  end
end


string linebuf568 = "";
logic hitMadPrint568 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc568_inst_done && ((spc568_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint568 = 1;
       linebuf568 = {linebuf568, spc568_phy_pc_w[8:1]};
       if (spc568_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 568, linebuf568);
          linebuf568 = "";
       end
    end else begin
       hitMadPrint568 = 0;
    end
  end
end


string linebuf569 = "";
logic hitMadPrint569 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc569_inst_done && ((spc569_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint569 = 1;
       linebuf569 = {linebuf569, spc569_phy_pc_w[8:1]};
       if (spc569_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 569, linebuf569);
          linebuf569 = "";
       end
    end else begin
       hitMadPrint569 = 0;
    end
  end
end


string linebuf570 = "";
logic hitMadPrint570 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc570_inst_done && ((spc570_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint570 = 1;
       linebuf570 = {linebuf570, spc570_phy_pc_w[8:1]};
       if (spc570_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 570, linebuf570);
          linebuf570 = "";
       end
    end else begin
       hitMadPrint570 = 0;
    end
  end
end


string linebuf571 = "";
logic hitMadPrint571 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc571_inst_done && ((spc571_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint571 = 1;
       linebuf571 = {linebuf571, spc571_phy_pc_w[8:1]};
       if (spc571_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 571, linebuf571);
          linebuf571 = "";
       end
    end else begin
       hitMadPrint571 = 0;
    end
  end
end


string linebuf572 = "";
logic hitMadPrint572 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc572_inst_done && ((spc572_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint572 = 1;
       linebuf572 = {linebuf572, spc572_phy_pc_w[8:1]};
       if (spc572_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 572, linebuf572);
          linebuf572 = "";
       end
    end else begin
       hitMadPrint572 = 0;
    end
  end
end


string linebuf573 = "";
logic hitMadPrint573 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc573_inst_done && ((spc573_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint573 = 1;
       linebuf573 = {linebuf573, spc573_phy_pc_w[8:1]};
       if (spc573_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 573, linebuf573);
          linebuf573 = "";
       end
    end else begin
       hitMadPrint573 = 0;
    end
  end
end


string linebuf574 = "";
logic hitMadPrint574 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc574_inst_done && ((spc574_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint574 = 1;
       linebuf574 = {linebuf574, spc574_phy_pc_w[8:1]};
       if (spc574_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 574, linebuf574);
          linebuf574 = "";
       end
    end else begin
       hitMadPrint574 = 0;
    end
  end
end


string linebuf575 = "";
logic hitMadPrint575 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc575_inst_done && ((spc575_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint575 = 1;
       linebuf575 = {linebuf575, spc575_phy_pc_w[8:1]};
       if (spc575_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 575, linebuf575);
          linebuf575 = "";
       end
    end else begin
       hitMadPrint575 = 0;
    end
  end
end


string linebuf576 = "";
logic hitMadPrint576 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc576_inst_done && ((spc576_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint576 = 1;
       linebuf576 = {linebuf576, spc576_phy_pc_w[8:1]};
       if (spc576_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 576, linebuf576);
          linebuf576 = "";
       end
    end else begin
       hitMadPrint576 = 0;
    end
  end
end


string linebuf577 = "";
logic hitMadPrint577 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc577_inst_done && ((spc577_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint577 = 1;
       linebuf577 = {linebuf577, spc577_phy_pc_w[8:1]};
       if (spc577_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 577, linebuf577);
          linebuf577 = "";
       end
    end else begin
       hitMadPrint577 = 0;
    end
  end
end


string linebuf578 = "";
logic hitMadPrint578 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc578_inst_done && ((spc578_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint578 = 1;
       linebuf578 = {linebuf578, spc578_phy_pc_w[8:1]};
       if (spc578_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 578, linebuf578);
          linebuf578 = "";
       end
    end else begin
       hitMadPrint578 = 0;
    end
  end
end


string linebuf579 = "";
logic hitMadPrint579 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc579_inst_done && ((spc579_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint579 = 1;
       linebuf579 = {linebuf579, spc579_phy_pc_w[8:1]};
       if (spc579_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 579, linebuf579);
          linebuf579 = "";
       end
    end else begin
       hitMadPrint579 = 0;
    end
  end
end


string linebuf580 = "";
logic hitMadPrint580 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc580_inst_done && ((spc580_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint580 = 1;
       linebuf580 = {linebuf580, spc580_phy_pc_w[8:1]};
       if (spc580_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 580, linebuf580);
          linebuf580 = "";
       end
    end else begin
       hitMadPrint580 = 0;
    end
  end
end


string linebuf581 = "";
logic hitMadPrint581 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc581_inst_done && ((spc581_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint581 = 1;
       linebuf581 = {linebuf581, spc581_phy_pc_w[8:1]};
       if (spc581_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 581, linebuf581);
          linebuf581 = "";
       end
    end else begin
       hitMadPrint581 = 0;
    end
  end
end


string linebuf582 = "";
logic hitMadPrint582 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc582_inst_done && ((spc582_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint582 = 1;
       linebuf582 = {linebuf582, spc582_phy_pc_w[8:1]};
       if (spc582_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 582, linebuf582);
          linebuf582 = "";
       end
    end else begin
       hitMadPrint582 = 0;
    end
  end
end


string linebuf583 = "";
logic hitMadPrint583 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc583_inst_done && ((spc583_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint583 = 1;
       linebuf583 = {linebuf583, spc583_phy_pc_w[8:1]};
       if (spc583_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 583, linebuf583);
          linebuf583 = "";
       end
    end else begin
       hitMadPrint583 = 0;
    end
  end
end


string linebuf584 = "";
logic hitMadPrint584 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc584_inst_done && ((spc584_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint584 = 1;
       linebuf584 = {linebuf584, spc584_phy_pc_w[8:1]};
       if (spc584_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 584, linebuf584);
          linebuf584 = "";
       end
    end else begin
       hitMadPrint584 = 0;
    end
  end
end


string linebuf585 = "";
logic hitMadPrint585 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc585_inst_done && ((spc585_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint585 = 1;
       linebuf585 = {linebuf585, spc585_phy_pc_w[8:1]};
       if (spc585_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 585, linebuf585);
          linebuf585 = "";
       end
    end else begin
       hitMadPrint585 = 0;
    end
  end
end


string linebuf586 = "";
logic hitMadPrint586 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc586_inst_done && ((spc586_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint586 = 1;
       linebuf586 = {linebuf586, spc586_phy_pc_w[8:1]};
       if (spc586_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 586, linebuf586);
          linebuf586 = "";
       end
    end else begin
       hitMadPrint586 = 0;
    end
  end
end


string linebuf587 = "";
logic hitMadPrint587 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc587_inst_done && ((spc587_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint587 = 1;
       linebuf587 = {linebuf587, spc587_phy_pc_w[8:1]};
       if (spc587_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 587, linebuf587);
          linebuf587 = "";
       end
    end else begin
       hitMadPrint587 = 0;
    end
  end
end


string linebuf588 = "";
logic hitMadPrint588 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc588_inst_done && ((spc588_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint588 = 1;
       linebuf588 = {linebuf588, spc588_phy_pc_w[8:1]};
       if (spc588_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 588, linebuf588);
          linebuf588 = "";
       end
    end else begin
       hitMadPrint588 = 0;
    end
  end
end


string linebuf589 = "";
logic hitMadPrint589 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc589_inst_done && ((spc589_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint589 = 1;
       linebuf589 = {linebuf589, spc589_phy_pc_w[8:1]};
       if (spc589_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 589, linebuf589);
          linebuf589 = "";
       end
    end else begin
       hitMadPrint589 = 0;
    end
  end
end


string linebuf590 = "";
logic hitMadPrint590 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc590_inst_done && ((spc590_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint590 = 1;
       linebuf590 = {linebuf590, spc590_phy_pc_w[8:1]};
       if (spc590_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 590, linebuf590);
          linebuf590 = "";
       end
    end else begin
       hitMadPrint590 = 0;
    end
  end
end


string linebuf591 = "";
logic hitMadPrint591 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc591_inst_done && ((spc591_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint591 = 1;
       linebuf591 = {linebuf591, spc591_phy_pc_w[8:1]};
       if (spc591_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 591, linebuf591);
          linebuf591 = "";
       end
    end else begin
       hitMadPrint591 = 0;
    end
  end
end


string linebuf592 = "";
logic hitMadPrint592 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc592_inst_done && ((spc592_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint592 = 1;
       linebuf592 = {linebuf592, spc592_phy_pc_w[8:1]};
       if (spc592_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 592, linebuf592);
          linebuf592 = "";
       end
    end else begin
       hitMadPrint592 = 0;
    end
  end
end


string linebuf593 = "";
logic hitMadPrint593 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc593_inst_done && ((spc593_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint593 = 1;
       linebuf593 = {linebuf593, spc593_phy_pc_w[8:1]};
       if (spc593_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 593, linebuf593);
          linebuf593 = "";
       end
    end else begin
       hitMadPrint593 = 0;
    end
  end
end


string linebuf594 = "";
logic hitMadPrint594 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc594_inst_done && ((spc594_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint594 = 1;
       linebuf594 = {linebuf594, spc594_phy_pc_w[8:1]};
       if (spc594_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 594, linebuf594);
          linebuf594 = "";
       end
    end else begin
       hitMadPrint594 = 0;
    end
  end
end


string linebuf595 = "";
logic hitMadPrint595 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc595_inst_done && ((spc595_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint595 = 1;
       linebuf595 = {linebuf595, spc595_phy_pc_w[8:1]};
       if (spc595_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 595, linebuf595);
          linebuf595 = "";
       end
    end else begin
       hitMadPrint595 = 0;
    end
  end
end


string linebuf596 = "";
logic hitMadPrint596 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc596_inst_done && ((spc596_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint596 = 1;
       linebuf596 = {linebuf596, spc596_phy_pc_w[8:1]};
       if (spc596_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 596, linebuf596);
          linebuf596 = "";
       end
    end else begin
       hitMadPrint596 = 0;
    end
  end
end


string linebuf597 = "";
logic hitMadPrint597 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc597_inst_done && ((spc597_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint597 = 1;
       linebuf597 = {linebuf597, spc597_phy_pc_w[8:1]};
       if (spc597_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 597, linebuf597);
          linebuf597 = "";
       end
    end else begin
       hitMadPrint597 = 0;
    end
  end
end


string linebuf598 = "";
logic hitMadPrint598 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc598_inst_done && ((spc598_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint598 = 1;
       linebuf598 = {linebuf598, spc598_phy_pc_w[8:1]};
       if (spc598_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 598, linebuf598);
          linebuf598 = "";
       end
    end else begin
       hitMadPrint598 = 0;
    end
  end
end


string linebuf599 = "";
logic hitMadPrint599 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc599_inst_done && ((spc599_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint599 = 1;
       linebuf599 = {linebuf599, spc599_phy_pc_w[8:1]};
       if (spc599_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 599, linebuf599);
          linebuf599 = "";
       end
    end else begin
       hitMadPrint599 = 0;
    end
  end
end


string linebuf600 = "";
logic hitMadPrint600 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc600_inst_done && ((spc600_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint600 = 1;
       linebuf600 = {linebuf600, spc600_phy_pc_w[8:1]};
       if (spc600_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 600, linebuf600);
          linebuf600 = "";
       end
    end else begin
       hitMadPrint600 = 0;
    end
  end
end


string linebuf601 = "";
logic hitMadPrint601 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc601_inst_done && ((spc601_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint601 = 1;
       linebuf601 = {linebuf601, spc601_phy_pc_w[8:1]};
       if (spc601_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 601, linebuf601);
          linebuf601 = "";
       end
    end else begin
       hitMadPrint601 = 0;
    end
  end
end


string linebuf602 = "";
logic hitMadPrint602 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc602_inst_done && ((spc602_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint602 = 1;
       linebuf602 = {linebuf602, spc602_phy_pc_w[8:1]};
       if (spc602_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 602, linebuf602);
          linebuf602 = "";
       end
    end else begin
       hitMadPrint602 = 0;
    end
  end
end


string linebuf603 = "";
logic hitMadPrint603 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc603_inst_done && ((spc603_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint603 = 1;
       linebuf603 = {linebuf603, spc603_phy_pc_w[8:1]};
       if (spc603_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 603, linebuf603);
          linebuf603 = "";
       end
    end else begin
       hitMadPrint603 = 0;
    end
  end
end


string linebuf604 = "";
logic hitMadPrint604 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc604_inst_done && ((spc604_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint604 = 1;
       linebuf604 = {linebuf604, spc604_phy_pc_w[8:1]};
       if (spc604_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 604, linebuf604);
          linebuf604 = "";
       end
    end else begin
       hitMadPrint604 = 0;
    end
  end
end


string linebuf605 = "";
logic hitMadPrint605 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc605_inst_done && ((spc605_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint605 = 1;
       linebuf605 = {linebuf605, spc605_phy_pc_w[8:1]};
       if (spc605_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 605, linebuf605);
          linebuf605 = "";
       end
    end else begin
       hitMadPrint605 = 0;
    end
  end
end


string linebuf606 = "";
logic hitMadPrint606 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc606_inst_done && ((spc606_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint606 = 1;
       linebuf606 = {linebuf606, spc606_phy_pc_w[8:1]};
       if (spc606_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 606, linebuf606);
          linebuf606 = "";
       end
    end else begin
       hitMadPrint606 = 0;
    end
  end
end


string linebuf607 = "";
logic hitMadPrint607 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc607_inst_done && ((spc607_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint607 = 1;
       linebuf607 = {linebuf607, spc607_phy_pc_w[8:1]};
       if (spc607_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 607, linebuf607);
          linebuf607 = "";
       end
    end else begin
       hitMadPrint607 = 0;
    end
  end
end


string linebuf608 = "";
logic hitMadPrint608 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc608_inst_done && ((spc608_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint608 = 1;
       linebuf608 = {linebuf608, spc608_phy_pc_w[8:1]};
       if (spc608_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 608, linebuf608);
          linebuf608 = "";
       end
    end else begin
       hitMadPrint608 = 0;
    end
  end
end


string linebuf609 = "";
logic hitMadPrint609 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc609_inst_done && ((spc609_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint609 = 1;
       linebuf609 = {linebuf609, spc609_phy_pc_w[8:1]};
       if (spc609_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 609, linebuf609);
          linebuf609 = "";
       end
    end else begin
       hitMadPrint609 = 0;
    end
  end
end


string linebuf610 = "";
logic hitMadPrint610 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc610_inst_done && ((spc610_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint610 = 1;
       linebuf610 = {linebuf610, spc610_phy_pc_w[8:1]};
       if (spc610_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 610, linebuf610);
          linebuf610 = "";
       end
    end else begin
       hitMadPrint610 = 0;
    end
  end
end


string linebuf611 = "";
logic hitMadPrint611 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc611_inst_done && ((spc611_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint611 = 1;
       linebuf611 = {linebuf611, spc611_phy_pc_w[8:1]};
       if (spc611_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 611, linebuf611);
          linebuf611 = "";
       end
    end else begin
       hitMadPrint611 = 0;
    end
  end
end


string linebuf612 = "";
logic hitMadPrint612 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc612_inst_done && ((spc612_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint612 = 1;
       linebuf612 = {linebuf612, spc612_phy_pc_w[8:1]};
       if (spc612_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 612, linebuf612);
          linebuf612 = "";
       end
    end else begin
       hitMadPrint612 = 0;
    end
  end
end


string linebuf613 = "";
logic hitMadPrint613 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc613_inst_done && ((spc613_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint613 = 1;
       linebuf613 = {linebuf613, spc613_phy_pc_w[8:1]};
       if (spc613_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 613, linebuf613);
          linebuf613 = "";
       end
    end else begin
       hitMadPrint613 = 0;
    end
  end
end


string linebuf614 = "";
logic hitMadPrint614 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc614_inst_done && ((spc614_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint614 = 1;
       linebuf614 = {linebuf614, spc614_phy_pc_w[8:1]};
       if (spc614_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 614, linebuf614);
          linebuf614 = "";
       end
    end else begin
       hitMadPrint614 = 0;
    end
  end
end


string linebuf615 = "";
logic hitMadPrint615 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc615_inst_done && ((spc615_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint615 = 1;
       linebuf615 = {linebuf615, spc615_phy_pc_w[8:1]};
       if (spc615_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 615, linebuf615);
          linebuf615 = "";
       end
    end else begin
       hitMadPrint615 = 0;
    end
  end
end


string linebuf616 = "";
logic hitMadPrint616 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc616_inst_done && ((spc616_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint616 = 1;
       linebuf616 = {linebuf616, spc616_phy_pc_w[8:1]};
       if (spc616_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 616, linebuf616);
          linebuf616 = "";
       end
    end else begin
       hitMadPrint616 = 0;
    end
  end
end


string linebuf617 = "";
logic hitMadPrint617 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc617_inst_done && ((spc617_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint617 = 1;
       linebuf617 = {linebuf617, spc617_phy_pc_w[8:1]};
       if (spc617_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 617, linebuf617);
          linebuf617 = "";
       end
    end else begin
       hitMadPrint617 = 0;
    end
  end
end


string linebuf618 = "";
logic hitMadPrint618 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc618_inst_done && ((spc618_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint618 = 1;
       linebuf618 = {linebuf618, spc618_phy_pc_w[8:1]};
       if (spc618_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 618, linebuf618);
          linebuf618 = "";
       end
    end else begin
       hitMadPrint618 = 0;
    end
  end
end


string linebuf619 = "";
logic hitMadPrint619 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc619_inst_done && ((spc619_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint619 = 1;
       linebuf619 = {linebuf619, spc619_phy_pc_w[8:1]};
       if (spc619_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 619, linebuf619);
          linebuf619 = "";
       end
    end else begin
       hitMadPrint619 = 0;
    end
  end
end


string linebuf620 = "";
logic hitMadPrint620 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc620_inst_done && ((spc620_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint620 = 1;
       linebuf620 = {linebuf620, spc620_phy_pc_w[8:1]};
       if (spc620_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 620, linebuf620);
          linebuf620 = "";
       end
    end else begin
       hitMadPrint620 = 0;
    end
  end
end


string linebuf621 = "";
logic hitMadPrint621 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc621_inst_done && ((spc621_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint621 = 1;
       linebuf621 = {linebuf621, spc621_phy_pc_w[8:1]};
       if (spc621_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 621, linebuf621);
          linebuf621 = "";
       end
    end else begin
       hitMadPrint621 = 0;
    end
  end
end


string linebuf622 = "";
logic hitMadPrint622 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc622_inst_done && ((spc622_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint622 = 1;
       linebuf622 = {linebuf622, spc622_phy_pc_w[8:1]};
       if (spc622_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 622, linebuf622);
          linebuf622 = "";
       end
    end else begin
       hitMadPrint622 = 0;
    end
  end
end


string linebuf623 = "";
logic hitMadPrint623 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc623_inst_done && ((spc623_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint623 = 1;
       linebuf623 = {linebuf623, spc623_phy_pc_w[8:1]};
       if (spc623_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 623, linebuf623);
          linebuf623 = "";
       end
    end else begin
       hitMadPrint623 = 0;
    end
  end
end


string linebuf624 = "";
logic hitMadPrint624 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc624_inst_done && ((spc624_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint624 = 1;
       linebuf624 = {linebuf624, spc624_phy_pc_w[8:1]};
       if (spc624_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 624, linebuf624);
          linebuf624 = "";
       end
    end else begin
       hitMadPrint624 = 0;
    end
  end
end


string linebuf625 = "";
logic hitMadPrint625 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc625_inst_done && ((spc625_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint625 = 1;
       linebuf625 = {linebuf625, spc625_phy_pc_w[8:1]};
       if (spc625_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 625, linebuf625);
          linebuf625 = "";
       end
    end else begin
       hitMadPrint625 = 0;
    end
  end
end


string linebuf626 = "";
logic hitMadPrint626 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc626_inst_done && ((spc626_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint626 = 1;
       linebuf626 = {linebuf626, spc626_phy_pc_w[8:1]};
       if (spc626_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 626, linebuf626);
          linebuf626 = "";
       end
    end else begin
       hitMadPrint626 = 0;
    end
  end
end


string linebuf627 = "";
logic hitMadPrint627 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc627_inst_done && ((spc627_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint627 = 1;
       linebuf627 = {linebuf627, spc627_phy_pc_w[8:1]};
       if (spc627_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 627, linebuf627);
          linebuf627 = "";
       end
    end else begin
       hitMadPrint627 = 0;
    end
  end
end


string linebuf628 = "";
logic hitMadPrint628 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc628_inst_done && ((spc628_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint628 = 1;
       linebuf628 = {linebuf628, spc628_phy_pc_w[8:1]};
       if (spc628_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 628, linebuf628);
          linebuf628 = "";
       end
    end else begin
       hitMadPrint628 = 0;
    end
  end
end


string linebuf629 = "";
logic hitMadPrint629 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc629_inst_done && ((spc629_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint629 = 1;
       linebuf629 = {linebuf629, spc629_phy_pc_w[8:1]};
       if (spc629_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 629, linebuf629);
          linebuf629 = "";
       end
    end else begin
       hitMadPrint629 = 0;
    end
  end
end


string linebuf630 = "";
logic hitMadPrint630 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc630_inst_done && ((spc630_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint630 = 1;
       linebuf630 = {linebuf630, spc630_phy_pc_w[8:1]};
       if (spc630_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 630, linebuf630);
          linebuf630 = "";
       end
    end else begin
       hitMadPrint630 = 0;
    end
  end
end


string linebuf631 = "";
logic hitMadPrint631 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc631_inst_done && ((spc631_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint631 = 1;
       linebuf631 = {linebuf631, spc631_phy_pc_w[8:1]};
       if (spc631_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 631, linebuf631);
          linebuf631 = "";
       end
    end else begin
       hitMadPrint631 = 0;
    end
  end
end


string linebuf632 = "";
logic hitMadPrint632 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc632_inst_done && ((spc632_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint632 = 1;
       linebuf632 = {linebuf632, spc632_phy_pc_w[8:1]};
       if (spc632_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 632, linebuf632);
          linebuf632 = "";
       end
    end else begin
       hitMadPrint632 = 0;
    end
  end
end


string linebuf633 = "";
logic hitMadPrint633 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc633_inst_done && ((spc633_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint633 = 1;
       linebuf633 = {linebuf633, spc633_phy_pc_w[8:1]};
       if (spc633_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 633, linebuf633);
          linebuf633 = "";
       end
    end else begin
       hitMadPrint633 = 0;
    end
  end
end


string linebuf634 = "";
logic hitMadPrint634 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc634_inst_done && ((spc634_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint634 = 1;
       linebuf634 = {linebuf634, spc634_phy_pc_w[8:1]};
       if (spc634_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 634, linebuf634);
          linebuf634 = "";
       end
    end else begin
       hitMadPrint634 = 0;
    end
  end
end


string linebuf635 = "";
logic hitMadPrint635 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc635_inst_done && ((spc635_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint635 = 1;
       linebuf635 = {linebuf635, spc635_phy_pc_w[8:1]};
       if (spc635_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 635, linebuf635);
          linebuf635 = "";
       end
    end else begin
       hitMadPrint635 = 0;
    end
  end
end


string linebuf636 = "";
logic hitMadPrint636 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc636_inst_done && ((spc636_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint636 = 1;
       linebuf636 = {linebuf636, spc636_phy_pc_w[8:1]};
       if (spc636_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 636, linebuf636);
          linebuf636 = "";
       end
    end else begin
       hitMadPrint636 = 0;
    end
  end
end


string linebuf637 = "";
logic hitMadPrint637 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc637_inst_done && ((spc637_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint637 = 1;
       linebuf637 = {linebuf637, spc637_phy_pc_w[8:1]};
       if (spc637_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 637, linebuf637);
          linebuf637 = "";
       end
    end else begin
       hitMadPrint637 = 0;
    end
  end
end


string linebuf638 = "";
logic hitMadPrint638 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc638_inst_done && ((spc638_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint638 = 1;
       linebuf638 = {linebuf638, spc638_phy_pc_w[8:1]};
       if (spc638_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 638, linebuf638);
          linebuf638 = "";
       end
    end else begin
       hitMadPrint638 = 0;
    end
  end
end


string linebuf639 = "";
logic hitMadPrint639 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc639_inst_done && ((spc639_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint639 = 1;
       linebuf639 = {linebuf639, spc639_phy_pc_w[8:1]};
       if (spc639_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 639, linebuf639);
          linebuf639 = "";
       end
    end else begin
       hitMadPrint639 = 0;
    end
  end
end


string linebuf640 = "";
logic hitMadPrint640 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc640_inst_done && ((spc640_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint640 = 1;
       linebuf640 = {linebuf640, spc640_phy_pc_w[8:1]};
       if (spc640_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 640, linebuf640);
          linebuf640 = "";
       end
    end else begin
       hitMadPrint640 = 0;
    end
  end
end


string linebuf641 = "";
logic hitMadPrint641 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc641_inst_done && ((spc641_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint641 = 1;
       linebuf641 = {linebuf641, spc641_phy_pc_w[8:1]};
       if (spc641_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 641, linebuf641);
          linebuf641 = "";
       end
    end else begin
       hitMadPrint641 = 0;
    end
  end
end


string linebuf642 = "";
logic hitMadPrint642 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc642_inst_done && ((spc642_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint642 = 1;
       linebuf642 = {linebuf642, spc642_phy_pc_w[8:1]};
       if (spc642_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 642, linebuf642);
          linebuf642 = "";
       end
    end else begin
       hitMadPrint642 = 0;
    end
  end
end


string linebuf643 = "";
logic hitMadPrint643 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc643_inst_done && ((spc643_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint643 = 1;
       linebuf643 = {linebuf643, spc643_phy_pc_w[8:1]};
       if (spc643_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 643, linebuf643);
          linebuf643 = "";
       end
    end else begin
       hitMadPrint643 = 0;
    end
  end
end


string linebuf644 = "";
logic hitMadPrint644 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc644_inst_done && ((spc644_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint644 = 1;
       linebuf644 = {linebuf644, spc644_phy_pc_w[8:1]};
       if (spc644_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 644, linebuf644);
          linebuf644 = "";
       end
    end else begin
       hitMadPrint644 = 0;
    end
  end
end


string linebuf645 = "";
logic hitMadPrint645 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc645_inst_done && ((spc645_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint645 = 1;
       linebuf645 = {linebuf645, spc645_phy_pc_w[8:1]};
       if (spc645_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 645, linebuf645);
          linebuf645 = "";
       end
    end else begin
       hitMadPrint645 = 0;
    end
  end
end


string linebuf646 = "";
logic hitMadPrint646 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc646_inst_done && ((spc646_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint646 = 1;
       linebuf646 = {linebuf646, spc646_phy_pc_w[8:1]};
       if (spc646_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 646, linebuf646);
          linebuf646 = "";
       end
    end else begin
       hitMadPrint646 = 0;
    end
  end
end


string linebuf647 = "";
logic hitMadPrint647 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc647_inst_done && ((spc647_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint647 = 1;
       linebuf647 = {linebuf647, spc647_phy_pc_w[8:1]};
       if (spc647_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 647, linebuf647);
          linebuf647 = "";
       end
    end else begin
       hitMadPrint647 = 0;
    end
  end
end


string linebuf648 = "";
logic hitMadPrint648 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc648_inst_done && ((spc648_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint648 = 1;
       linebuf648 = {linebuf648, spc648_phy_pc_w[8:1]};
       if (spc648_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 648, linebuf648);
          linebuf648 = "";
       end
    end else begin
       hitMadPrint648 = 0;
    end
  end
end


string linebuf649 = "";
logic hitMadPrint649 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc649_inst_done && ((spc649_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint649 = 1;
       linebuf649 = {linebuf649, spc649_phy_pc_w[8:1]};
       if (spc649_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 649, linebuf649);
          linebuf649 = "";
       end
    end else begin
       hitMadPrint649 = 0;
    end
  end
end


string linebuf650 = "";
logic hitMadPrint650 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc650_inst_done && ((spc650_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint650 = 1;
       linebuf650 = {linebuf650, spc650_phy_pc_w[8:1]};
       if (spc650_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 650, linebuf650);
          linebuf650 = "";
       end
    end else begin
       hitMadPrint650 = 0;
    end
  end
end


string linebuf651 = "";
logic hitMadPrint651 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc651_inst_done && ((spc651_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint651 = 1;
       linebuf651 = {linebuf651, spc651_phy_pc_w[8:1]};
       if (spc651_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 651, linebuf651);
          linebuf651 = "";
       end
    end else begin
       hitMadPrint651 = 0;
    end
  end
end


string linebuf652 = "";
logic hitMadPrint652 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc652_inst_done && ((spc652_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint652 = 1;
       linebuf652 = {linebuf652, spc652_phy_pc_w[8:1]};
       if (spc652_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 652, linebuf652);
          linebuf652 = "";
       end
    end else begin
       hitMadPrint652 = 0;
    end
  end
end


string linebuf653 = "";
logic hitMadPrint653 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc653_inst_done && ((spc653_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint653 = 1;
       linebuf653 = {linebuf653, spc653_phy_pc_w[8:1]};
       if (spc653_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 653, linebuf653);
          linebuf653 = "";
       end
    end else begin
       hitMadPrint653 = 0;
    end
  end
end


string linebuf654 = "";
logic hitMadPrint654 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc654_inst_done && ((spc654_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint654 = 1;
       linebuf654 = {linebuf654, spc654_phy_pc_w[8:1]};
       if (spc654_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 654, linebuf654);
          linebuf654 = "";
       end
    end else begin
       hitMadPrint654 = 0;
    end
  end
end


string linebuf655 = "";
logic hitMadPrint655 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc655_inst_done && ((spc655_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint655 = 1;
       linebuf655 = {linebuf655, spc655_phy_pc_w[8:1]};
       if (spc655_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 655, linebuf655);
          linebuf655 = "";
       end
    end else begin
       hitMadPrint655 = 0;
    end
  end
end


string linebuf656 = "";
logic hitMadPrint656 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc656_inst_done && ((spc656_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint656 = 1;
       linebuf656 = {linebuf656, spc656_phy_pc_w[8:1]};
       if (spc656_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 656, linebuf656);
          linebuf656 = "";
       end
    end else begin
       hitMadPrint656 = 0;
    end
  end
end


string linebuf657 = "";
logic hitMadPrint657 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc657_inst_done && ((spc657_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint657 = 1;
       linebuf657 = {linebuf657, spc657_phy_pc_w[8:1]};
       if (spc657_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 657, linebuf657);
          linebuf657 = "";
       end
    end else begin
       hitMadPrint657 = 0;
    end
  end
end


string linebuf658 = "";
logic hitMadPrint658 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc658_inst_done && ((spc658_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint658 = 1;
       linebuf658 = {linebuf658, spc658_phy_pc_w[8:1]};
       if (spc658_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 658, linebuf658);
          linebuf658 = "";
       end
    end else begin
       hitMadPrint658 = 0;
    end
  end
end


string linebuf659 = "";
logic hitMadPrint659 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc659_inst_done && ((spc659_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint659 = 1;
       linebuf659 = {linebuf659, spc659_phy_pc_w[8:1]};
       if (spc659_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 659, linebuf659);
          linebuf659 = "";
       end
    end else begin
       hitMadPrint659 = 0;
    end
  end
end


string linebuf660 = "";
logic hitMadPrint660 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc660_inst_done && ((spc660_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint660 = 1;
       linebuf660 = {linebuf660, spc660_phy_pc_w[8:1]};
       if (spc660_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 660, linebuf660);
          linebuf660 = "";
       end
    end else begin
       hitMadPrint660 = 0;
    end
  end
end


string linebuf661 = "";
logic hitMadPrint661 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc661_inst_done && ((spc661_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint661 = 1;
       linebuf661 = {linebuf661, spc661_phy_pc_w[8:1]};
       if (spc661_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 661, linebuf661);
          linebuf661 = "";
       end
    end else begin
       hitMadPrint661 = 0;
    end
  end
end


string linebuf662 = "";
logic hitMadPrint662 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc662_inst_done && ((spc662_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint662 = 1;
       linebuf662 = {linebuf662, spc662_phy_pc_w[8:1]};
       if (spc662_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 662, linebuf662);
          linebuf662 = "";
       end
    end else begin
       hitMadPrint662 = 0;
    end
  end
end


string linebuf663 = "";
logic hitMadPrint663 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc663_inst_done && ((spc663_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint663 = 1;
       linebuf663 = {linebuf663, spc663_phy_pc_w[8:1]};
       if (spc663_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 663, linebuf663);
          linebuf663 = "";
       end
    end else begin
       hitMadPrint663 = 0;
    end
  end
end


string linebuf664 = "";
logic hitMadPrint664 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc664_inst_done && ((spc664_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint664 = 1;
       linebuf664 = {linebuf664, spc664_phy_pc_w[8:1]};
       if (spc664_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 664, linebuf664);
          linebuf664 = "";
       end
    end else begin
       hitMadPrint664 = 0;
    end
  end
end


string linebuf665 = "";
logic hitMadPrint665 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc665_inst_done && ((spc665_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint665 = 1;
       linebuf665 = {linebuf665, spc665_phy_pc_w[8:1]};
       if (spc665_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 665, linebuf665);
          linebuf665 = "";
       end
    end else begin
       hitMadPrint665 = 0;
    end
  end
end


string linebuf666 = "";
logic hitMadPrint666 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc666_inst_done && ((spc666_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint666 = 1;
       linebuf666 = {linebuf666, spc666_phy_pc_w[8:1]};
       if (spc666_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 666, linebuf666);
          linebuf666 = "";
       end
    end else begin
       hitMadPrint666 = 0;
    end
  end
end


string linebuf667 = "";
logic hitMadPrint667 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc667_inst_done && ((spc667_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint667 = 1;
       linebuf667 = {linebuf667, spc667_phy_pc_w[8:1]};
       if (spc667_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 667, linebuf667);
          linebuf667 = "";
       end
    end else begin
       hitMadPrint667 = 0;
    end
  end
end


string linebuf668 = "";
logic hitMadPrint668 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc668_inst_done && ((spc668_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint668 = 1;
       linebuf668 = {linebuf668, spc668_phy_pc_w[8:1]};
       if (spc668_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 668, linebuf668);
          linebuf668 = "";
       end
    end else begin
       hitMadPrint668 = 0;
    end
  end
end


string linebuf669 = "";
logic hitMadPrint669 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc669_inst_done && ((spc669_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint669 = 1;
       linebuf669 = {linebuf669, spc669_phy_pc_w[8:1]};
       if (spc669_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 669, linebuf669);
          linebuf669 = "";
       end
    end else begin
       hitMadPrint669 = 0;
    end
  end
end


string linebuf670 = "";
logic hitMadPrint670 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc670_inst_done && ((spc670_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint670 = 1;
       linebuf670 = {linebuf670, spc670_phy_pc_w[8:1]};
       if (spc670_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 670, linebuf670);
          linebuf670 = "";
       end
    end else begin
       hitMadPrint670 = 0;
    end
  end
end


string linebuf671 = "";
logic hitMadPrint671 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc671_inst_done && ((spc671_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint671 = 1;
       linebuf671 = {linebuf671, spc671_phy_pc_w[8:1]};
       if (spc671_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 671, linebuf671);
          linebuf671 = "";
       end
    end else begin
       hitMadPrint671 = 0;
    end
  end
end


string linebuf672 = "";
logic hitMadPrint672 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc672_inst_done && ((spc672_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint672 = 1;
       linebuf672 = {linebuf672, spc672_phy_pc_w[8:1]};
       if (spc672_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 672, linebuf672);
          linebuf672 = "";
       end
    end else begin
       hitMadPrint672 = 0;
    end
  end
end


string linebuf673 = "";
logic hitMadPrint673 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc673_inst_done && ((spc673_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint673 = 1;
       linebuf673 = {linebuf673, spc673_phy_pc_w[8:1]};
       if (spc673_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 673, linebuf673);
          linebuf673 = "";
       end
    end else begin
       hitMadPrint673 = 0;
    end
  end
end


string linebuf674 = "";
logic hitMadPrint674 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc674_inst_done && ((spc674_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint674 = 1;
       linebuf674 = {linebuf674, spc674_phy_pc_w[8:1]};
       if (spc674_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 674, linebuf674);
          linebuf674 = "";
       end
    end else begin
       hitMadPrint674 = 0;
    end
  end
end


string linebuf675 = "";
logic hitMadPrint675 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc675_inst_done && ((spc675_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint675 = 1;
       linebuf675 = {linebuf675, spc675_phy_pc_w[8:1]};
       if (spc675_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 675, linebuf675);
          linebuf675 = "";
       end
    end else begin
       hitMadPrint675 = 0;
    end
  end
end


string linebuf676 = "";
logic hitMadPrint676 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc676_inst_done && ((spc676_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint676 = 1;
       linebuf676 = {linebuf676, spc676_phy_pc_w[8:1]};
       if (spc676_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 676, linebuf676);
          linebuf676 = "";
       end
    end else begin
       hitMadPrint676 = 0;
    end
  end
end


string linebuf677 = "";
logic hitMadPrint677 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc677_inst_done && ((spc677_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint677 = 1;
       linebuf677 = {linebuf677, spc677_phy_pc_w[8:1]};
       if (spc677_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 677, linebuf677);
          linebuf677 = "";
       end
    end else begin
       hitMadPrint677 = 0;
    end
  end
end


string linebuf678 = "";
logic hitMadPrint678 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc678_inst_done && ((spc678_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint678 = 1;
       linebuf678 = {linebuf678, spc678_phy_pc_w[8:1]};
       if (spc678_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 678, linebuf678);
          linebuf678 = "";
       end
    end else begin
       hitMadPrint678 = 0;
    end
  end
end


string linebuf679 = "";
logic hitMadPrint679 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc679_inst_done && ((spc679_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint679 = 1;
       linebuf679 = {linebuf679, spc679_phy_pc_w[8:1]};
       if (spc679_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 679, linebuf679);
          linebuf679 = "";
       end
    end else begin
       hitMadPrint679 = 0;
    end
  end
end


string linebuf680 = "";
logic hitMadPrint680 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc680_inst_done && ((spc680_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint680 = 1;
       linebuf680 = {linebuf680, spc680_phy_pc_w[8:1]};
       if (spc680_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 680, linebuf680);
          linebuf680 = "";
       end
    end else begin
       hitMadPrint680 = 0;
    end
  end
end


string linebuf681 = "";
logic hitMadPrint681 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc681_inst_done && ((spc681_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint681 = 1;
       linebuf681 = {linebuf681, spc681_phy_pc_w[8:1]};
       if (spc681_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 681, linebuf681);
          linebuf681 = "";
       end
    end else begin
       hitMadPrint681 = 0;
    end
  end
end


string linebuf682 = "";
logic hitMadPrint682 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc682_inst_done && ((spc682_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint682 = 1;
       linebuf682 = {linebuf682, spc682_phy_pc_w[8:1]};
       if (spc682_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 682, linebuf682);
          linebuf682 = "";
       end
    end else begin
       hitMadPrint682 = 0;
    end
  end
end


string linebuf683 = "";
logic hitMadPrint683 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc683_inst_done && ((spc683_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint683 = 1;
       linebuf683 = {linebuf683, spc683_phy_pc_w[8:1]};
       if (spc683_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 683, linebuf683);
          linebuf683 = "";
       end
    end else begin
       hitMadPrint683 = 0;
    end
  end
end


string linebuf684 = "";
logic hitMadPrint684 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc684_inst_done && ((spc684_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint684 = 1;
       linebuf684 = {linebuf684, spc684_phy_pc_w[8:1]};
       if (spc684_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 684, linebuf684);
          linebuf684 = "";
       end
    end else begin
       hitMadPrint684 = 0;
    end
  end
end


string linebuf685 = "";
logic hitMadPrint685 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc685_inst_done && ((spc685_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint685 = 1;
       linebuf685 = {linebuf685, spc685_phy_pc_w[8:1]};
       if (spc685_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 685, linebuf685);
          linebuf685 = "";
       end
    end else begin
       hitMadPrint685 = 0;
    end
  end
end


string linebuf686 = "";
logic hitMadPrint686 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc686_inst_done && ((spc686_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint686 = 1;
       linebuf686 = {linebuf686, spc686_phy_pc_w[8:1]};
       if (spc686_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 686, linebuf686);
          linebuf686 = "";
       end
    end else begin
       hitMadPrint686 = 0;
    end
  end
end


string linebuf687 = "";
logic hitMadPrint687 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc687_inst_done && ((spc687_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint687 = 1;
       linebuf687 = {linebuf687, spc687_phy_pc_w[8:1]};
       if (spc687_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 687, linebuf687);
          linebuf687 = "";
       end
    end else begin
       hitMadPrint687 = 0;
    end
  end
end


string linebuf688 = "";
logic hitMadPrint688 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc688_inst_done && ((spc688_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint688 = 1;
       linebuf688 = {linebuf688, spc688_phy_pc_w[8:1]};
       if (spc688_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 688, linebuf688);
          linebuf688 = "";
       end
    end else begin
       hitMadPrint688 = 0;
    end
  end
end


string linebuf689 = "";
logic hitMadPrint689 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc689_inst_done && ((spc689_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint689 = 1;
       linebuf689 = {linebuf689, spc689_phy_pc_w[8:1]};
       if (spc689_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 689, linebuf689);
          linebuf689 = "";
       end
    end else begin
       hitMadPrint689 = 0;
    end
  end
end


string linebuf690 = "";
logic hitMadPrint690 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc690_inst_done && ((spc690_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint690 = 1;
       linebuf690 = {linebuf690, spc690_phy_pc_w[8:1]};
       if (spc690_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 690, linebuf690);
          linebuf690 = "";
       end
    end else begin
       hitMadPrint690 = 0;
    end
  end
end


string linebuf691 = "";
logic hitMadPrint691 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc691_inst_done && ((spc691_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint691 = 1;
       linebuf691 = {linebuf691, spc691_phy_pc_w[8:1]};
       if (spc691_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 691, linebuf691);
          linebuf691 = "";
       end
    end else begin
       hitMadPrint691 = 0;
    end
  end
end


string linebuf692 = "";
logic hitMadPrint692 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc692_inst_done && ((spc692_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint692 = 1;
       linebuf692 = {linebuf692, spc692_phy_pc_w[8:1]};
       if (spc692_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 692, linebuf692);
          linebuf692 = "";
       end
    end else begin
       hitMadPrint692 = 0;
    end
  end
end


string linebuf693 = "";
logic hitMadPrint693 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc693_inst_done && ((spc693_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint693 = 1;
       linebuf693 = {linebuf693, spc693_phy_pc_w[8:1]};
       if (spc693_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 693, linebuf693);
          linebuf693 = "";
       end
    end else begin
       hitMadPrint693 = 0;
    end
  end
end


string linebuf694 = "";
logic hitMadPrint694 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc694_inst_done && ((spc694_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint694 = 1;
       linebuf694 = {linebuf694, spc694_phy_pc_w[8:1]};
       if (spc694_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 694, linebuf694);
          linebuf694 = "";
       end
    end else begin
       hitMadPrint694 = 0;
    end
  end
end


string linebuf695 = "";
logic hitMadPrint695 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc695_inst_done && ((spc695_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint695 = 1;
       linebuf695 = {linebuf695, spc695_phy_pc_w[8:1]};
       if (spc695_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 695, linebuf695);
          linebuf695 = "";
       end
    end else begin
       hitMadPrint695 = 0;
    end
  end
end


string linebuf696 = "";
logic hitMadPrint696 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc696_inst_done && ((spc696_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint696 = 1;
       linebuf696 = {linebuf696, spc696_phy_pc_w[8:1]};
       if (spc696_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 696, linebuf696);
          linebuf696 = "";
       end
    end else begin
       hitMadPrint696 = 0;
    end
  end
end


string linebuf697 = "";
logic hitMadPrint697 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc697_inst_done && ((spc697_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint697 = 1;
       linebuf697 = {linebuf697, spc697_phy_pc_w[8:1]};
       if (spc697_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 697, linebuf697);
          linebuf697 = "";
       end
    end else begin
       hitMadPrint697 = 0;
    end
  end
end


string linebuf698 = "";
logic hitMadPrint698 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc698_inst_done && ((spc698_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint698 = 1;
       linebuf698 = {linebuf698, spc698_phy_pc_w[8:1]};
       if (spc698_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 698, linebuf698);
          linebuf698 = "";
       end
    end else begin
       hitMadPrint698 = 0;
    end
  end
end


string linebuf699 = "";
logic hitMadPrint699 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc699_inst_done && ((spc699_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint699 = 1;
       linebuf699 = {linebuf699, spc699_phy_pc_w[8:1]};
       if (spc699_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 699, linebuf699);
          linebuf699 = "";
       end
    end else begin
       hitMadPrint699 = 0;
    end
  end
end


string linebuf700 = "";
logic hitMadPrint700 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc700_inst_done && ((spc700_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint700 = 1;
       linebuf700 = {linebuf700, spc700_phy_pc_w[8:1]};
       if (spc700_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 700, linebuf700);
          linebuf700 = "";
       end
    end else begin
       hitMadPrint700 = 0;
    end
  end
end


string linebuf701 = "";
logic hitMadPrint701 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc701_inst_done && ((spc701_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint701 = 1;
       linebuf701 = {linebuf701, spc701_phy_pc_w[8:1]};
       if (spc701_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 701, linebuf701);
          linebuf701 = "";
       end
    end else begin
       hitMadPrint701 = 0;
    end
  end
end


string linebuf702 = "";
logic hitMadPrint702 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc702_inst_done && ((spc702_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint702 = 1;
       linebuf702 = {linebuf702, spc702_phy_pc_w[8:1]};
       if (spc702_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 702, linebuf702);
          linebuf702 = "";
       end
    end else begin
       hitMadPrint702 = 0;
    end
  end
end


string linebuf703 = "";
logic hitMadPrint703 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc703_inst_done && ((spc703_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint703 = 1;
       linebuf703 = {linebuf703, spc703_phy_pc_w[8:1]};
       if (spc703_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 703, linebuf703);
          linebuf703 = "";
       end
    end else begin
       hitMadPrint703 = 0;
    end
  end
end


string linebuf704 = "";
logic hitMadPrint704 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc704_inst_done && ((spc704_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint704 = 1;
       linebuf704 = {linebuf704, spc704_phy_pc_w[8:1]};
       if (spc704_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 704, linebuf704);
          linebuf704 = "";
       end
    end else begin
       hitMadPrint704 = 0;
    end
  end
end


string linebuf705 = "";
logic hitMadPrint705 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc705_inst_done && ((spc705_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint705 = 1;
       linebuf705 = {linebuf705, spc705_phy_pc_w[8:1]};
       if (spc705_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 705, linebuf705);
          linebuf705 = "";
       end
    end else begin
       hitMadPrint705 = 0;
    end
  end
end


string linebuf706 = "";
logic hitMadPrint706 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc706_inst_done && ((spc706_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint706 = 1;
       linebuf706 = {linebuf706, spc706_phy_pc_w[8:1]};
       if (spc706_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 706, linebuf706);
          linebuf706 = "";
       end
    end else begin
       hitMadPrint706 = 0;
    end
  end
end


string linebuf707 = "";
logic hitMadPrint707 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc707_inst_done && ((spc707_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint707 = 1;
       linebuf707 = {linebuf707, spc707_phy_pc_w[8:1]};
       if (spc707_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 707, linebuf707);
          linebuf707 = "";
       end
    end else begin
       hitMadPrint707 = 0;
    end
  end
end


string linebuf708 = "";
logic hitMadPrint708 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc708_inst_done && ((spc708_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint708 = 1;
       linebuf708 = {linebuf708, spc708_phy_pc_w[8:1]};
       if (spc708_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 708, linebuf708);
          linebuf708 = "";
       end
    end else begin
       hitMadPrint708 = 0;
    end
  end
end


string linebuf709 = "";
logic hitMadPrint709 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc709_inst_done && ((spc709_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint709 = 1;
       linebuf709 = {linebuf709, spc709_phy_pc_w[8:1]};
       if (spc709_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 709, linebuf709);
          linebuf709 = "";
       end
    end else begin
       hitMadPrint709 = 0;
    end
  end
end


string linebuf710 = "";
logic hitMadPrint710 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc710_inst_done && ((spc710_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint710 = 1;
       linebuf710 = {linebuf710, spc710_phy_pc_w[8:1]};
       if (spc710_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 710, linebuf710);
          linebuf710 = "";
       end
    end else begin
       hitMadPrint710 = 0;
    end
  end
end


string linebuf711 = "";
logic hitMadPrint711 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc711_inst_done && ((spc711_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint711 = 1;
       linebuf711 = {linebuf711, spc711_phy_pc_w[8:1]};
       if (spc711_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 711, linebuf711);
          linebuf711 = "";
       end
    end else begin
       hitMadPrint711 = 0;
    end
  end
end


string linebuf712 = "";
logic hitMadPrint712 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc712_inst_done && ((spc712_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint712 = 1;
       linebuf712 = {linebuf712, spc712_phy_pc_w[8:1]};
       if (spc712_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 712, linebuf712);
          linebuf712 = "";
       end
    end else begin
       hitMadPrint712 = 0;
    end
  end
end


string linebuf713 = "";
logic hitMadPrint713 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc713_inst_done && ((spc713_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint713 = 1;
       linebuf713 = {linebuf713, spc713_phy_pc_w[8:1]};
       if (spc713_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 713, linebuf713);
          linebuf713 = "";
       end
    end else begin
       hitMadPrint713 = 0;
    end
  end
end


string linebuf714 = "";
logic hitMadPrint714 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc714_inst_done && ((spc714_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint714 = 1;
       linebuf714 = {linebuf714, spc714_phy_pc_w[8:1]};
       if (spc714_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 714, linebuf714);
          linebuf714 = "";
       end
    end else begin
       hitMadPrint714 = 0;
    end
  end
end


string linebuf715 = "";
logic hitMadPrint715 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc715_inst_done && ((spc715_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint715 = 1;
       linebuf715 = {linebuf715, spc715_phy_pc_w[8:1]};
       if (spc715_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 715, linebuf715);
          linebuf715 = "";
       end
    end else begin
       hitMadPrint715 = 0;
    end
  end
end


string linebuf716 = "";
logic hitMadPrint716 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc716_inst_done && ((spc716_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint716 = 1;
       linebuf716 = {linebuf716, spc716_phy_pc_w[8:1]};
       if (spc716_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 716, linebuf716);
          linebuf716 = "";
       end
    end else begin
       hitMadPrint716 = 0;
    end
  end
end


string linebuf717 = "";
logic hitMadPrint717 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc717_inst_done && ((spc717_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint717 = 1;
       linebuf717 = {linebuf717, spc717_phy_pc_w[8:1]};
       if (spc717_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 717, linebuf717);
          linebuf717 = "";
       end
    end else begin
       hitMadPrint717 = 0;
    end
  end
end


string linebuf718 = "";
logic hitMadPrint718 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc718_inst_done && ((spc718_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint718 = 1;
       linebuf718 = {linebuf718, spc718_phy_pc_w[8:1]};
       if (spc718_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 718, linebuf718);
          linebuf718 = "";
       end
    end else begin
       hitMadPrint718 = 0;
    end
  end
end


string linebuf719 = "";
logic hitMadPrint719 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc719_inst_done && ((spc719_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint719 = 1;
       linebuf719 = {linebuf719, spc719_phy_pc_w[8:1]};
       if (spc719_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 719, linebuf719);
          linebuf719 = "";
       end
    end else begin
       hitMadPrint719 = 0;
    end
  end
end


string linebuf720 = "";
logic hitMadPrint720 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc720_inst_done && ((spc720_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint720 = 1;
       linebuf720 = {linebuf720, spc720_phy_pc_w[8:1]};
       if (spc720_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 720, linebuf720);
          linebuf720 = "";
       end
    end else begin
       hitMadPrint720 = 0;
    end
  end
end


string linebuf721 = "";
logic hitMadPrint721 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc721_inst_done && ((spc721_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint721 = 1;
       linebuf721 = {linebuf721, spc721_phy_pc_w[8:1]};
       if (spc721_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 721, linebuf721);
          linebuf721 = "";
       end
    end else begin
       hitMadPrint721 = 0;
    end
  end
end


string linebuf722 = "";
logic hitMadPrint722 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc722_inst_done && ((spc722_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint722 = 1;
       linebuf722 = {linebuf722, spc722_phy_pc_w[8:1]};
       if (spc722_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 722, linebuf722);
          linebuf722 = "";
       end
    end else begin
       hitMadPrint722 = 0;
    end
  end
end


string linebuf723 = "";
logic hitMadPrint723 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc723_inst_done && ((spc723_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint723 = 1;
       linebuf723 = {linebuf723, spc723_phy_pc_w[8:1]};
       if (spc723_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 723, linebuf723);
          linebuf723 = "";
       end
    end else begin
       hitMadPrint723 = 0;
    end
  end
end


string linebuf724 = "";
logic hitMadPrint724 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc724_inst_done && ((spc724_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint724 = 1;
       linebuf724 = {linebuf724, spc724_phy_pc_w[8:1]};
       if (spc724_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 724, linebuf724);
          linebuf724 = "";
       end
    end else begin
       hitMadPrint724 = 0;
    end
  end
end


string linebuf725 = "";
logic hitMadPrint725 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc725_inst_done && ((spc725_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint725 = 1;
       linebuf725 = {linebuf725, spc725_phy_pc_w[8:1]};
       if (spc725_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 725, linebuf725);
          linebuf725 = "";
       end
    end else begin
       hitMadPrint725 = 0;
    end
  end
end


string linebuf726 = "";
logic hitMadPrint726 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc726_inst_done && ((spc726_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint726 = 1;
       linebuf726 = {linebuf726, spc726_phy_pc_w[8:1]};
       if (spc726_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 726, linebuf726);
          linebuf726 = "";
       end
    end else begin
       hitMadPrint726 = 0;
    end
  end
end


string linebuf727 = "";
logic hitMadPrint727 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc727_inst_done && ((spc727_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint727 = 1;
       linebuf727 = {linebuf727, spc727_phy_pc_w[8:1]};
       if (spc727_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 727, linebuf727);
          linebuf727 = "";
       end
    end else begin
       hitMadPrint727 = 0;
    end
  end
end


string linebuf728 = "";
logic hitMadPrint728 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc728_inst_done && ((spc728_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint728 = 1;
       linebuf728 = {linebuf728, spc728_phy_pc_w[8:1]};
       if (spc728_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 728, linebuf728);
          linebuf728 = "";
       end
    end else begin
       hitMadPrint728 = 0;
    end
  end
end


string linebuf729 = "";
logic hitMadPrint729 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc729_inst_done && ((spc729_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint729 = 1;
       linebuf729 = {linebuf729, spc729_phy_pc_w[8:1]};
       if (spc729_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 729, linebuf729);
          linebuf729 = "";
       end
    end else begin
       hitMadPrint729 = 0;
    end
  end
end


string linebuf730 = "";
logic hitMadPrint730 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc730_inst_done && ((spc730_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint730 = 1;
       linebuf730 = {linebuf730, spc730_phy_pc_w[8:1]};
       if (spc730_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 730, linebuf730);
          linebuf730 = "";
       end
    end else begin
       hitMadPrint730 = 0;
    end
  end
end


string linebuf731 = "";
logic hitMadPrint731 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc731_inst_done && ((spc731_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint731 = 1;
       linebuf731 = {linebuf731, spc731_phy_pc_w[8:1]};
       if (spc731_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 731, linebuf731);
          linebuf731 = "";
       end
    end else begin
       hitMadPrint731 = 0;
    end
  end
end


string linebuf732 = "";
logic hitMadPrint732 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc732_inst_done && ((spc732_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint732 = 1;
       linebuf732 = {linebuf732, spc732_phy_pc_w[8:1]};
       if (spc732_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 732, linebuf732);
          linebuf732 = "";
       end
    end else begin
       hitMadPrint732 = 0;
    end
  end
end


string linebuf733 = "";
logic hitMadPrint733 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc733_inst_done && ((spc733_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint733 = 1;
       linebuf733 = {linebuf733, spc733_phy_pc_w[8:1]};
       if (spc733_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 733, linebuf733);
          linebuf733 = "";
       end
    end else begin
       hitMadPrint733 = 0;
    end
  end
end


string linebuf734 = "";
logic hitMadPrint734 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc734_inst_done && ((spc734_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint734 = 1;
       linebuf734 = {linebuf734, spc734_phy_pc_w[8:1]};
       if (spc734_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 734, linebuf734);
          linebuf734 = "";
       end
    end else begin
       hitMadPrint734 = 0;
    end
  end
end


string linebuf735 = "";
logic hitMadPrint735 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc735_inst_done && ((spc735_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint735 = 1;
       linebuf735 = {linebuf735, spc735_phy_pc_w[8:1]};
       if (spc735_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 735, linebuf735);
          linebuf735 = "";
       end
    end else begin
       hitMadPrint735 = 0;
    end
  end
end


string linebuf736 = "";
logic hitMadPrint736 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc736_inst_done && ((spc736_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint736 = 1;
       linebuf736 = {linebuf736, spc736_phy_pc_w[8:1]};
       if (spc736_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 736, linebuf736);
          linebuf736 = "";
       end
    end else begin
       hitMadPrint736 = 0;
    end
  end
end


string linebuf737 = "";
logic hitMadPrint737 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc737_inst_done && ((spc737_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint737 = 1;
       linebuf737 = {linebuf737, spc737_phy_pc_w[8:1]};
       if (spc737_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 737, linebuf737);
          linebuf737 = "";
       end
    end else begin
       hitMadPrint737 = 0;
    end
  end
end


string linebuf738 = "";
logic hitMadPrint738 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc738_inst_done && ((spc738_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint738 = 1;
       linebuf738 = {linebuf738, spc738_phy_pc_w[8:1]};
       if (spc738_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 738, linebuf738);
          linebuf738 = "";
       end
    end else begin
       hitMadPrint738 = 0;
    end
  end
end


string linebuf739 = "";
logic hitMadPrint739 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc739_inst_done && ((spc739_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint739 = 1;
       linebuf739 = {linebuf739, spc739_phy_pc_w[8:1]};
       if (spc739_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 739, linebuf739);
          linebuf739 = "";
       end
    end else begin
       hitMadPrint739 = 0;
    end
  end
end


string linebuf740 = "";
logic hitMadPrint740 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc740_inst_done && ((spc740_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint740 = 1;
       linebuf740 = {linebuf740, spc740_phy_pc_w[8:1]};
       if (spc740_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 740, linebuf740);
          linebuf740 = "";
       end
    end else begin
       hitMadPrint740 = 0;
    end
  end
end


string linebuf741 = "";
logic hitMadPrint741 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc741_inst_done && ((spc741_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint741 = 1;
       linebuf741 = {linebuf741, spc741_phy_pc_w[8:1]};
       if (spc741_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 741, linebuf741);
          linebuf741 = "";
       end
    end else begin
       hitMadPrint741 = 0;
    end
  end
end


string linebuf742 = "";
logic hitMadPrint742 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc742_inst_done && ((spc742_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint742 = 1;
       linebuf742 = {linebuf742, spc742_phy_pc_w[8:1]};
       if (spc742_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 742, linebuf742);
          linebuf742 = "";
       end
    end else begin
       hitMadPrint742 = 0;
    end
  end
end


string linebuf743 = "";
logic hitMadPrint743 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc743_inst_done && ((spc743_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint743 = 1;
       linebuf743 = {linebuf743, spc743_phy_pc_w[8:1]};
       if (spc743_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 743, linebuf743);
          linebuf743 = "";
       end
    end else begin
       hitMadPrint743 = 0;
    end
  end
end


string linebuf744 = "";
logic hitMadPrint744 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc744_inst_done && ((spc744_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint744 = 1;
       linebuf744 = {linebuf744, spc744_phy_pc_w[8:1]};
       if (spc744_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 744, linebuf744);
          linebuf744 = "";
       end
    end else begin
       hitMadPrint744 = 0;
    end
  end
end


string linebuf745 = "";
logic hitMadPrint745 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc745_inst_done && ((spc745_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint745 = 1;
       linebuf745 = {linebuf745, spc745_phy_pc_w[8:1]};
       if (spc745_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 745, linebuf745);
          linebuf745 = "";
       end
    end else begin
       hitMadPrint745 = 0;
    end
  end
end


string linebuf746 = "";
logic hitMadPrint746 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc746_inst_done && ((spc746_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint746 = 1;
       linebuf746 = {linebuf746, spc746_phy_pc_w[8:1]};
       if (spc746_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 746, linebuf746);
          linebuf746 = "";
       end
    end else begin
       hitMadPrint746 = 0;
    end
  end
end


string linebuf747 = "";
logic hitMadPrint747 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc747_inst_done && ((spc747_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint747 = 1;
       linebuf747 = {linebuf747, spc747_phy_pc_w[8:1]};
       if (spc747_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 747, linebuf747);
          linebuf747 = "";
       end
    end else begin
       hitMadPrint747 = 0;
    end
  end
end


string linebuf748 = "";
logic hitMadPrint748 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc748_inst_done && ((spc748_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint748 = 1;
       linebuf748 = {linebuf748, spc748_phy_pc_w[8:1]};
       if (spc748_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 748, linebuf748);
          linebuf748 = "";
       end
    end else begin
       hitMadPrint748 = 0;
    end
  end
end


string linebuf749 = "";
logic hitMadPrint749 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc749_inst_done && ((spc749_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint749 = 1;
       linebuf749 = {linebuf749, spc749_phy_pc_w[8:1]};
       if (spc749_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 749, linebuf749);
          linebuf749 = "";
       end
    end else begin
       hitMadPrint749 = 0;
    end
  end
end


string linebuf750 = "";
logic hitMadPrint750 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc750_inst_done && ((spc750_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint750 = 1;
       linebuf750 = {linebuf750, spc750_phy_pc_w[8:1]};
       if (spc750_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 750, linebuf750);
          linebuf750 = "";
       end
    end else begin
       hitMadPrint750 = 0;
    end
  end
end


string linebuf751 = "";
logic hitMadPrint751 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc751_inst_done && ((spc751_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint751 = 1;
       linebuf751 = {linebuf751, spc751_phy_pc_w[8:1]};
       if (spc751_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 751, linebuf751);
          linebuf751 = "";
       end
    end else begin
       hitMadPrint751 = 0;
    end
  end
end


string linebuf752 = "";
logic hitMadPrint752 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc752_inst_done && ((spc752_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint752 = 1;
       linebuf752 = {linebuf752, spc752_phy_pc_w[8:1]};
       if (spc752_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 752, linebuf752);
          linebuf752 = "";
       end
    end else begin
       hitMadPrint752 = 0;
    end
  end
end


string linebuf753 = "";
logic hitMadPrint753 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc753_inst_done && ((spc753_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint753 = 1;
       linebuf753 = {linebuf753, spc753_phy_pc_w[8:1]};
       if (spc753_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 753, linebuf753);
          linebuf753 = "";
       end
    end else begin
       hitMadPrint753 = 0;
    end
  end
end


string linebuf754 = "";
logic hitMadPrint754 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc754_inst_done && ((spc754_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint754 = 1;
       linebuf754 = {linebuf754, spc754_phy_pc_w[8:1]};
       if (spc754_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 754, linebuf754);
          linebuf754 = "";
       end
    end else begin
       hitMadPrint754 = 0;
    end
  end
end


string linebuf755 = "";
logic hitMadPrint755 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc755_inst_done && ((spc755_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint755 = 1;
       linebuf755 = {linebuf755, spc755_phy_pc_w[8:1]};
       if (spc755_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 755, linebuf755);
          linebuf755 = "";
       end
    end else begin
       hitMadPrint755 = 0;
    end
  end
end


string linebuf756 = "";
logic hitMadPrint756 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc756_inst_done && ((spc756_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint756 = 1;
       linebuf756 = {linebuf756, spc756_phy_pc_w[8:1]};
       if (spc756_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 756, linebuf756);
          linebuf756 = "";
       end
    end else begin
       hitMadPrint756 = 0;
    end
  end
end


string linebuf757 = "";
logic hitMadPrint757 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc757_inst_done && ((spc757_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint757 = 1;
       linebuf757 = {linebuf757, spc757_phy_pc_w[8:1]};
       if (spc757_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 757, linebuf757);
          linebuf757 = "";
       end
    end else begin
       hitMadPrint757 = 0;
    end
  end
end


string linebuf758 = "";
logic hitMadPrint758 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc758_inst_done && ((spc758_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint758 = 1;
       linebuf758 = {linebuf758, spc758_phy_pc_w[8:1]};
       if (spc758_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 758, linebuf758);
          linebuf758 = "";
       end
    end else begin
       hitMadPrint758 = 0;
    end
  end
end


string linebuf759 = "";
logic hitMadPrint759 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc759_inst_done && ((spc759_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint759 = 1;
       linebuf759 = {linebuf759, spc759_phy_pc_w[8:1]};
       if (spc759_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 759, linebuf759);
          linebuf759 = "";
       end
    end else begin
       hitMadPrint759 = 0;
    end
  end
end


string linebuf760 = "";
logic hitMadPrint760 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc760_inst_done && ((spc760_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint760 = 1;
       linebuf760 = {linebuf760, spc760_phy_pc_w[8:1]};
       if (spc760_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 760, linebuf760);
          linebuf760 = "";
       end
    end else begin
       hitMadPrint760 = 0;
    end
  end
end


string linebuf761 = "";
logic hitMadPrint761 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc761_inst_done && ((spc761_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint761 = 1;
       linebuf761 = {linebuf761, spc761_phy_pc_w[8:1]};
       if (spc761_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 761, linebuf761);
          linebuf761 = "";
       end
    end else begin
       hitMadPrint761 = 0;
    end
  end
end


string linebuf762 = "";
logic hitMadPrint762 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc762_inst_done && ((spc762_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint762 = 1;
       linebuf762 = {linebuf762, spc762_phy_pc_w[8:1]};
       if (spc762_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 762, linebuf762);
          linebuf762 = "";
       end
    end else begin
       hitMadPrint762 = 0;
    end
  end
end


string linebuf763 = "";
logic hitMadPrint763 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc763_inst_done && ((spc763_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint763 = 1;
       linebuf763 = {linebuf763, spc763_phy_pc_w[8:1]};
       if (spc763_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 763, linebuf763);
          linebuf763 = "";
       end
    end else begin
       hitMadPrint763 = 0;
    end
  end
end


string linebuf764 = "";
logic hitMadPrint764 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc764_inst_done && ((spc764_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint764 = 1;
       linebuf764 = {linebuf764, spc764_phy_pc_w[8:1]};
       if (spc764_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 764, linebuf764);
          linebuf764 = "";
       end
    end else begin
       hitMadPrint764 = 0;
    end
  end
end


string linebuf765 = "";
logic hitMadPrint765 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc765_inst_done && ((spc765_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint765 = 1;
       linebuf765 = {linebuf765, spc765_phy_pc_w[8:1]};
       if (spc765_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 765, linebuf765);
          linebuf765 = "";
       end
    end else begin
       hitMadPrint765 = 0;
    end
  end
end


string linebuf766 = "";
logic hitMadPrint766 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc766_inst_done && ((spc766_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint766 = 1;
       linebuf766 = {linebuf766, spc766_phy_pc_w[8:1]};
       if (spc766_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 766, linebuf766);
          linebuf766 = "";
       end
    end else begin
       hitMadPrint766 = 0;
    end
  end
end


string linebuf767 = "";
logic hitMadPrint767 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc767_inst_done && ((spc767_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint767 = 1;
       linebuf767 = {linebuf767, spc767_phy_pc_w[8:1]};
       if (spc767_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 767, linebuf767);
          linebuf767 = "";
       end
    end else begin
       hitMadPrint767 = 0;
    end
  end
end


string linebuf768 = "";
logic hitMadPrint768 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc768_inst_done && ((spc768_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint768 = 1;
       linebuf768 = {linebuf768, spc768_phy_pc_w[8:1]};
       if (spc768_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 768, linebuf768);
          linebuf768 = "";
       end
    end else begin
       hitMadPrint768 = 0;
    end
  end
end


string linebuf769 = "";
logic hitMadPrint769 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc769_inst_done && ((spc769_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint769 = 1;
       linebuf769 = {linebuf769, spc769_phy_pc_w[8:1]};
       if (spc769_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 769, linebuf769);
          linebuf769 = "";
       end
    end else begin
       hitMadPrint769 = 0;
    end
  end
end


string linebuf770 = "";
logic hitMadPrint770 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc770_inst_done && ((spc770_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint770 = 1;
       linebuf770 = {linebuf770, spc770_phy_pc_w[8:1]};
       if (spc770_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 770, linebuf770);
          linebuf770 = "";
       end
    end else begin
       hitMadPrint770 = 0;
    end
  end
end


string linebuf771 = "";
logic hitMadPrint771 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc771_inst_done && ((spc771_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint771 = 1;
       linebuf771 = {linebuf771, spc771_phy_pc_w[8:1]};
       if (spc771_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 771, linebuf771);
          linebuf771 = "";
       end
    end else begin
       hitMadPrint771 = 0;
    end
  end
end


string linebuf772 = "";
logic hitMadPrint772 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc772_inst_done && ((spc772_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint772 = 1;
       linebuf772 = {linebuf772, spc772_phy_pc_w[8:1]};
       if (spc772_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 772, linebuf772);
          linebuf772 = "";
       end
    end else begin
       hitMadPrint772 = 0;
    end
  end
end


string linebuf773 = "";
logic hitMadPrint773 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc773_inst_done && ((spc773_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint773 = 1;
       linebuf773 = {linebuf773, spc773_phy_pc_w[8:1]};
       if (spc773_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 773, linebuf773);
          linebuf773 = "";
       end
    end else begin
       hitMadPrint773 = 0;
    end
  end
end


string linebuf774 = "";
logic hitMadPrint774 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc774_inst_done && ((spc774_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint774 = 1;
       linebuf774 = {linebuf774, spc774_phy_pc_w[8:1]};
       if (spc774_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 774, linebuf774);
          linebuf774 = "";
       end
    end else begin
       hitMadPrint774 = 0;
    end
  end
end


string linebuf775 = "";
logic hitMadPrint775 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc775_inst_done && ((spc775_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint775 = 1;
       linebuf775 = {linebuf775, spc775_phy_pc_w[8:1]};
       if (spc775_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 775, linebuf775);
          linebuf775 = "";
       end
    end else begin
       hitMadPrint775 = 0;
    end
  end
end


string linebuf776 = "";
logic hitMadPrint776 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc776_inst_done && ((spc776_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint776 = 1;
       linebuf776 = {linebuf776, spc776_phy_pc_w[8:1]};
       if (spc776_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 776, linebuf776);
          linebuf776 = "";
       end
    end else begin
       hitMadPrint776 = 0;
    end
  end
end


string linebuf777 = "";
logic hitMadPrint777 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc777_inst_done && ((spc777_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint777 = 1;
       linebuf777 = {linebuf777, spc777_phy_pc_w[8:1]};
       if (spc777_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 777, linebuf777);
          linebuf777 = "";
       end
    end else begin
       hitMadPrint777 = 0;
    end
  end
end


string linebuf778 = "";
logic hitMadPrint778 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc778_inst_done && ((spc778_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint778 = 1;
       linebuf778 = {linebuf778, spc778_phy_pc_w[8:1]};
       if (spc778_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 778, linebuf778);
          linebuf778 = "";
       end
    end else begin
       hitMadPrint778 = 0;
    end
  end
end


string linebuf779 = "";
logic hitMadPrint779 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc779_inst_done && ((spc779_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint779 = 1;
       linebuf779 = {linebuf779, spc779_phy_pc_w[8:1]};
       if (spc779_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 779, linebuf779);
          linebuf779 = "";
       end
    end else begin
       hitMadPrint779 = 0;
    end
  end
end


string linebuf780 = "";
logic hitMadPrint780 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc780_inst_done && ((spc780_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint780 = 1;
       linebuf780 = {linebuf780, spc780_phy_pc_w[8:1]};
       if (spc780_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 780, linebuf780);
          linebuf780 = "";
       end
    end else begin
       hitMadPrint780 = 0;
    end
  end
end


string linebuf781 = "";
logic hitMadPrint781 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc781_inst_done && ((spc781_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint781 = 1;
       linebuf781 = {linebuf781, spc781_phy_pc_w[8:1]};
       if (spc781_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 781, linebuf781);
          linebuf781 = "";
       end
    end else begin
       hitMadPrint781 = 0;
    end
  end
end


string linebuf782 = "";
logic hitMadPrint782 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc782_inst_done && ((spc782_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint782 = 1;
       linebuf782 = {linebuf782, spc782_phy_pc_w[8:1]};
       if (spc782_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 782, linebuf782);
          linebuf782 = "";
       end
    end else begin
       hitMadPrint782 = 0;
    end
  end
end


string linebuf783 = "";
logic hitMadPrint783 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc783_inst_done && ((spc783_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint783 = 1;
       linebuf783 = {linebuf783, spc783_phy_pc_w[8:1]};
       if (spc783_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 783, linebuf783);
          linebuf783 = "";
       end
    end else begin
       hitMadPrint783 = 0;
    end
  end
end


string linebuf784 = "";
logic hitMadPrint784 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc784_inst_done && ((spc784_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint784 = 1;
       linebuf784 = {linebuf784, spc784_phy_pc_w[8:1]};
       if (spc784_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 784, linebuf784);
          linebuf784 = "";
       end
    end else begin
       hitMadPrint784 = 0;
    end
  end
end


string linebuf785 = "";
logic hitMadPrint785 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc785_inst_done && ((spc785_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint785 = 1;
       linebuf785 = {linebuf785, spc785_phy_pc_w[8:1]};
       if (spc785_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 785, linebuf785);
          linebuf785 = "";
       end
    end else begin
       hitMadPrint785 = 0;
    end
  end
end


string linebuf786 = "";
logic hitMadPrint786 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc786_inst_done && ((spc786_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint786 = 1;
       linebuf786 = {linebuf786, spc786_phy_pc_w[8:1]};
       if (spc786_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 786, linebuf786);
          linebuf786 = "";
       end
    end else begin
       hitMadPrint786 = 0;
    end
  end
end


string linebuf787 = "";
logic hitMadPrint787 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc787_inst_done && ((spc787_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint787 = 1;
       linebuf787 = {linebuf787, spc787_phy_pc_w[8:1]};
       if (spc787_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 787, linebuf787);
          linebuf787 = "";
       end
    end else begin
       hitMadPrint787 = 0;
    end
  end
end


string linebuf788 = "";
logic hitMadPrint788 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc788_inst_done && ((spc788_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint788 = 1;
       linebuf788 = {linebuf788, spc788_phy_pc_w[8:1]};
       if (spc788_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 788, linebuf788);
          linebuf788 = "";
       end
    end else begin
       hitMadPrint788 = 0;
    end
  end
end


string linebuf789 = "";
logic hitMadPrint789 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc789_inst_done && ((spc789_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint789 = 1;
       linebuf789 = {linebuf789, spc789_phy_pc_w[8:1]};
       if (spc789_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 789, linebuf789);
          linebuf789 = "";
       end
    end else begin
       hitMadPrint789 = 0;
    end
  end
end


string linebuf790 = "";
logic hitMadPrint790 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc790_inst_done && ((spc790_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint790 = 1;
       linebuf790 = {linebuf790, spc790_phy_pc_w[8:1]};
       if (spc790_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 790, linebuf790);
          linebuf790 = "";
       end
    end else begin
       hitMadPrint790 = 0;
    end
  end
end


string linebuf791 = "";
logic hitMadPrint791 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc791_inst_done && ((spc791_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint791 = 1;
       linebuf791 = {linebuf791, spc791_phy_pc_w[8:1]};
       if (spc791_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 791, linebuf791);
          linebuf791 = "";
       end
    end else begin
       hitMadPrint791 = 0;
    end
  end
end


string linebuf792 = "";
logic hitMadPrint792 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc792_inst_done && ((spc792_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint792 = 1;
       linebuf792 = {linebuf792, spc792_phy_pc_w[8:1]};
       if (spc792_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 792, linebuf792);
          linebuf792 = "";
       end
    end else begin
       hitMadPrint792 = 0;
    end
  end
end


string linebuf793 = "";
logic hitMadPrint793 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc793_inst_done && ((spc793_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint793 = 1;
       linebuf793 = {linebuf793, spc793_phy_pc_w[8:1]};
       if (spc793_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 793, linebuf793);
          linebuf793 = "";
       end
    end else begin
       hitMadPrint793 = 0;
    end
  end
end


string linebuf794 = "";
logic hitMadPrint794 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc794_inst_done && ((spc794_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint794 = 1;
       linebuf794 = {linebuf794, spc794_phy_pc_w[8:1]};
       if (spc794_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 794, linebuf794);
          linebuf794 = "";
       end
    end else begin
       hitMadPrint794 = 0;
    end
  end
end


string linebuf795 = "";
logic hitMadPrint795 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc795_inst_done && ((spc795_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint795 = 1;
       linebuf795 = {linebuf795, spc795_phy_pc_w[8:1]};
       if (spc795_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 795, linebuf795);
          linebuf795 = "";
       end
    end else begin
       hitMadPrint795 = 0;
    end
  end
end


string linebuf796 = "";
logic hitMadPrint796 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc796_inst_done && ((spc796_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint796 = 1;
       linebuf796 = {linebuf796, spc796_phy_pc_w[8:1]};
       if (spc796_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 796, linebuf796);
          linebuf796 = "";
       end
    end else begin
       hitMadPrint796 = 0;
    end
  end
end


string linebuf797 = "";
logic hitMadPrint797 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc797_inst_done && ((spc797_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint797 = 1;
       linebuf797 = {linebuf797, spc797_phy_pc_w[8:1]};
       if (spc797_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 797, linebuf797);
          linebuf797 = "";
       end
    end else begin
       hitMadPrint797 = 0;
    end
  end
end


string linebuf798 = "";
logic hitMadPrint798 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc798_inst_done && ((spc798_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint798 = 1;
       linebuf798 = {linebuf798, spc798_phy_pc_w[8:1]};
       if (spc798_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 798, linebuf798);
          linebuf798 = "";
       end
    end else begin
       hitMadPrint798 = 0;
    end
  end
end


string linebuf799 = "";
logic hitMadPrint799 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc799_inst_done && ((spc799_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint799 = 1;
       linebuf799 = {linebuf799, spc799_phy_pc_w[8:1]};
       if (spc799_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 799, linebuf799);
          linebuf799 = "";
       end
    end else begin
       hitMadPrint799 = 0;
    end
  end
end


string linebuf800 = "";
logic hitMadPrint800 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc800_inst_done && ((spc800_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint800 = 1;
       linebuf800 = {linebuf800, spc800_phy_pc_w[8:1]};
       if (spc800_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 800, linebuf800);
          linebuf800 = "";
       end
    end else begin
       hitMadPrint800 = 0;
    end
  end
end


string linebuf801 = "";
logic hitMadPrint801 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc801_inst_done && ((spc801_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint801 = 1;
       linebuf801 = {linebuf801, spc801_phy_pc_w[8:1]};
       if (spc801_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 801, linebuf801);
          linebuf801 = "";
       end
    end else begin
       hitMadPrint801 = 0;
    end
  end
end


string linebuf802 = "";
logic hitMadPrint802 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc802_inst_done && ((spc802_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint802 = 1;
       linebuf802 = {linebuf802, spc802_phy_pc_w[8:1]};
       if (spc802_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 802, linebuf802);
          linebuf802 = "";
       end
    end else begin
       hitMadPrint802 = 0;
    end
  end
end


string linebuf803 = "";
logic hitMadPrint803 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc803_inst_done && ((spc803_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint803 = 1;
       linebuf803 = {linebuf803, spc803_phy_pc_w[8:1]};
       if (spc803_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 803, linebuf803);
          linebuf803 = "";
       end
    end else begin
       hitMadPrint803 = 0;
    end
  end
end


string linebuf804 = "";
logic hitMadPrint804 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc804_inst_done && ((spc804_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint804 = 1;
       linebuf804 = {linebuf804, spc804_phy_pc_w[8:1]};
       if (spc804_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 804, linebuf804);
          linebuf804 = "";
       end
    end else begin
       hitMadPrint804 = 0;
    end
  end
end


string linebuf805 = "";
logic hitMadPrint805 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc805_inst_done && ((spc805_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint805 = 1;
       linebuf805 = {linebuf805, spc805_phy_pc_w[8:1]};
       if (spc805_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 805, linebuf805);
          linebuf805 = "";
       end
    end else begin
       hitMadPrint805 = 0;
    end
  end
end


string linebuf806 = "";
logic hitMadPrint806 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc806_inst_done && ((spc806_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint806 = 1;
       linebuf806 = {linebuf806, spc806_phy_pc_w[8:1]};
       if (spc806_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 806, linebuf806);
          linebuf806 = "";
       end
    end else begin
       hitMadPrint806 = 0;
    end
  end
end


string linebuf807 = "";
logic hitMadPrint807 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc807_inst_done && ((spc807_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint807 = 1;
       linebuf807 = {linebuf807, spc807_phy_pc_w[8:1]};
       if (spc807_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 807, linebuf807);
          linebuf807 = "";
       end
    end else begin
       hitMadPrint807 = 0;
    end
  end
end


string linebuf808 = "";
logic hitMadPrint808 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc808_inst_done && ((spc808_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint808 = 1;
       linebuf808 = {linebuf808, spc808_phy_pc_w[8:1]};
       if (spc808_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 808, linebuf808);
          linebuf808 = "";
       end
    end else begin
       hitMadPrint808 = 0;
    end
  end
end


string linebuf809 = "";
logic hitMadPrint809 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc809_inst_done && ((spc809_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint809 = 1;
       linebuf809 = {linebuf809, spc809_phy_pc_w[8:1]};
       if (spc809_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 809, linebuf809);
          linebuf809 = "";
       end
    end else begin
       hitMadPrint809 = 0;
    end
  end
end


string linebuf810 = "";
logic hitMadPrint810 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc810_inst_done && ((spc810_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint810 = 1;
       linebuf810 = {linebuf810, spc810_phy_pc_w[8:1]};
       if (spc810_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 810, linebuf810);
          linebuf810 = "";
       end
    end else begin
       hitMadPrint810 = 0;
    end
  end
end


string linebuf811 = "";
logic hitMadPrint811 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc811_inst_done && ((spc811_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint811 = 1;
       linebuf811 = {linebuf811, spc811_phy_pc_w[8:1]};
       if (spc811_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 811, linebuf811);
          linebuf811 = "";
       end
    end else begin
       hitMadPrint811 = 0;
    end
  end
end


string linebuf812 = "";
logic hitMadPrint812 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc812_inst_done && ((spc812_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint812 = 1;
       linebuf812 = {linebuf812, spc812_phy_pc_w[8:1]};
       if (spc812_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 812, linebuf812);
          linebuf812 = "";
       end
    end else begin
       hitMadPrint812 = 0;
    end
  end
end


string linebuf813 = "";
logic hitMadPrint813 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc813_inst_done && ((spc813_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint813 = 1;
       linebuf813 = {linebuf813, spc813_phy_pc_w[8:1]};
       if (spc813_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 813, linebuf813);
          linebuf813 = "";
       end
    end else begin
       hitMadPrint813 = 0;
    end
  end
end


string linebuf814 = "";
logic hitMadPrint814 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc814_inst_done && ((spc814_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint814 = 1;
       linebuf814 = {linebuf814, spc814_phy_pc_w[8:1]};
       if (spc814_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 814, linebuf814);
          linebuf814 = "";
       end
    end else begin
       hitMadPrint814 = 0;
    end
  end
end


string linebuf815 = "";
logic hitMadPrint815 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc815_inst_done && ((spc815_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint815 = 1;
       linebuf815 = {linebuf815, spc815_phy_pc_w[8:1]};
       if (spc815_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 815, linebuf815);
          linebuf815 = "";
       end
    end else begin
       hitMadPrint815 = 0;
    end
  end
end


string linebuf816 = "";
logic hitMadPrint816 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc816_inst_done && ((spc816_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint816 = 1;
       linebuf816 = {linebuf816, spc816_phy_pc_w[8:1]};
       if (spc816_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 816, linebuf816);
          linebuf816 = "";
       end
    end else begin
       hitMadPrint816 = 0;
    end
  end
end


string linebuf817 = "";
logic hitMadPrint817 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc817_inst_done && ((spc817_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint817 = 1;
       linebuf817 = {linebuf817, spc817_phy_pc_w[8:1]};
       if (spc817_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 817, linebuf817);
          linebuf817 = "";
       end
    end else begin
       hitMadPrint817 = 0;
    end
  end
end


string linebuf818 = "";
logic hitMadPrint818 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc818_inst_done && ((spc818_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint818 = 1;
       linebuf818 = {linebuf818, spc818_phy_pc_w[8:1]};
       if (spc818_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 818, linebuf818);
          linebuf818 = "";
       end
    end else begin
       hitMadPrint818 = 0;
    end
  end
end


string linebuf819 = "";
logic hitMadPrint819 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc819_inst_done && ((spc819_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint819 = 1;
       linebuf819 = {linebuf819, spc819_phy_pc_w[8:1]};
       if (spc819_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 819, linebuf819);
          linebuf819 = "";
       end
    end else begin
       hitMadPrint819 = 0;
    end
  end
end


string linebuf820 = "";
logic hitMadPrint820 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc820_inst_done && ((spc820_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint820 = 1;
       linebuf820 = {linebuf820, spc820_phy_pc_w[8:1]};
       if (spc820_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 820, linebuf820);
          linebuf820 = "";
       end
    end else begin
       hitMadPrint820 = 0;
    end
  end
end


string linebuf821 = "";
logic hitMadPrint821 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc821_inst_done && ((spc821_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint821 = 1;
       linebuf821 = {linebuf821, spc821_phy_pc_w[8:1]};
       if (spc821_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 821, linebuf821);
          linebuf821 = "";
       end
    end else begin
       hitMadPrint821 = 0;
    end
  end
end


string linebuf822 = "";
logic hitMadPrint822 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc822_inst_done && ((spc822_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint822 = 1;
       linebuf822 = {linebuf822, spc822_phy_pc_w[8:1]};
       if (spc822_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 822, linebuf822);
          linebuf822 = "";
       end
    end else begin
       hitMadPrint822 = 0;
    end
  end
end


string linebuf823 = "";
logic hitMadPrint823 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc823_inst_done && ((spc823_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint823 = 1;
       linebuf823 = {linebuf823, spc823_phy_pc_w[8:1]};
       if (spc823_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 823, linebuf823);
          linebuf823 = "";
       end
    end else begin
       hitMadPrint823 = 0;
    end
  end
end


string linebuf824 = "";
logic hitMadPrint824 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc824_inst_done && ((spc824_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint824 = 1;
       linebuf824 = {linebuf824, spc824_phy_pc_w[8:1]};
       if (spc824_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 824, linebuf824);
          linebuf824 = "";
       end
    end else begin
       hitMadPrint824 = 0;
    end
  end
end


string linebuf825 = "";
logic hitMadPrint825 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc825_inst_done && ((spc825_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint825 = 1;
       linebuf825 = {linebuf825, spc825_phy_pc_w[8:1]};
       if (spc825_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 825, linebuf825);
          linebuf825 = "";
       end
    end else begin
       hitMadPrint825 = 0;
    end
  end
end


string linebuf826 = "";
logic hitMadPrint826 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc826_inst_done && ((spc826_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint826 = 1;
       linebuf826 = {linebuf826, spc826_phy_pc_w[8:1]};
       if (spc826_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 826, linebuf826);
          linebuf826 = "";
       end
    end else begin
       hitMadPrint826 = 0;
    end
  end
end


string linebuf827 = "";
logic hitMadPrint827 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc827_inst_done && ((spc827_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint827 = 1;
       linebuf827 = {linebuf827, spc827_phy_pc_w[8:1]};
       if (spc827_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 827, linebuf827);
          linebuf827 = "";
       end
    end else begin
       hitMadPrint827 = 0;
    end
  end
end


string linebuf828 = "";
logic hitMadPrint828 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc828_inst_done && ((spc828_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint828 = 1;
       linebuf828 = {linebuf828, spc828_phy_pc_w[8:1]};
       if (spc828_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 828, linebuf828);
          linebuf828 = "";
       end
    end else begin
       hitMadPrint828 = 0;
    end
  end
end


string linebuf829 = "";
logic hitMadPrint829 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc829_inst_done && ((spc829_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint829 = 1;
       linebuf829 = {linebuf829, spc829_phy_pc_w[8:1]};
       if (spc829_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 829, linebuf829);
          linebuf829 = "";
       end
    end else begin
       hitMadPrint829 = 0;
    end
  end
end


string linebuf830 = "";
logic hitMadPrint830 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc830_inst_done && ((spc830_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint830 = 1;
       linebuf830 = {linebuf830, spc830_phy_pc_w[8:1]};
       if (spc830_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 830, linebuf830);
          linebuf830 = "";
       end
    end else begin
       hitMadPrint830 = 0;
    end
  end
end


string linebuf831 = "";
logic hitMadPrint831 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc831_inst_done && ((spc831_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint831 = 1;
       linebuf831 = {linebuf831, spc831_phy_pc_w[8:1]};
       if (spc831_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 831, linebuf831);
          linebuf831 = "";
       end
    end else begin
       hitMadPrint831 = 0;
    end
  end
end


string linebuf832 = "";
logic hitMadPrint832 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc832_inst_done && ((spc832_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint832 = 1;
       linebuf832 = {linebuf832, spc832_phy_pc_w[8:1]};
       if (spc832_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 832, linebuf832);
          linebuf832 = "";
       end
    end else begin
       hitMadPrint832 = 0;
    end
  end
end


string linebuf833 = "";
logic hitMadPrint833 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc833_inst_done && ((spc833_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint833 = 1;
       linebuf833 = {linebuf833, spc833_phy_pc_w[8:1]};
       if (spc833_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 833, linebuf833);
          linebuf833 = "";
       end
    end else begin
       hitMadPrint833 = 0;
    end
  end
end


string linebuf834 = "";
logic hitMadPrint834 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc834_inst_done && ((spc834_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint834 = 1;
       linebuf834 = {linebuf834, spc834_phy_pc_w[8:1]};
       if (spc834_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 834, linebuf834);
          linebuf834 = "";
       end
    end else begin
       hitMadPrint834 = 0;
    end
  end
end


string linebuf835 = "";
logic hitMadPrint835 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc835_inst_done && ((spc835_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint835 = 1;
       linebuf835 = {linebuf835, spc835_phy_pc_w[8:1]};
       if (spc835_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 835, linebuf835);
          linebuf835 = "";
       end
    end else begin
       hitMadPrint835 = 0;
    end
  end
end


string linebuf836 = "";
logic hitMadPrint836 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc836_inst_done && ((spc836_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint836 = 1;
       linebuf836 = {linebuf836, spc836_phy_pc_w[8:1]};
       if (spc836_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 836, linebuf836);
          linebuf836 = "";
       end
    end else begin
       hitMadPrint836 = 0;
    end
  end
end


string linebuf837 = "";
logic hitMadPrint837 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc837_inst_done && ((spc837_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint837 = 1;
       linebuf837 = {linebuf837, spc837_phy_pc_w[8:1]};
       if (spc837_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 837, linebuf837);
          linebuf837 = "";
       end
    end else begin
       hitMadPrint837 = 0;
    end
  end
end


string linebuf838 = "";
logic hitMadPrint838 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc838_inst_done && ((spc838_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint838 = 1;
       linebuf838 = {linebuf838, spc838_phy_pc_w[8:1]};
       if (spc838_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 838, linebuf838);
          linebuf838 = "";
       end
    end else begin
       hitMadPrint838 = 0;
    end
  end
end


string linebuf839 = "";
logic hitMadPrint839 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc839_inst_done && ((spc839_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint839 = 1;
       linebuf839 = {linebuf839, spc839_phy_pc_w[8:1]};
       if (spc839_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 839, linebuf839);
          linebuf839 = "";
       end
    end else begin
       hitMadPrint839 = 0;
    end
  end
end


string linebuf840 = "";
logic hitMadPrint840 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc840_inst_done && ((spc840_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint840 = 1;
       linebuf840 = {linebuf840, spc840_phy_pc_w[8:1]};
       if (spc840_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 840, linebuf840);
          linebuf840 = "";
       end
    end else begin
       hitMadPrint840 = 0;
    end
  end
end


string linebuf841 = "";
logic hitMadPrint841 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc841_inst_done && ((spc841_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint841 = 1;
       linebuf841 = {linebuf841, spc841_phy_pc_w[8:1]};
       if (spc841_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 841, linebuf841);
          linebuf841 = "";
       end
    end else begin
       hitMadPrint841 = 0;
    end
  end
end


string linebuf842 = "";
logic hitMadPrint842 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc842_inst_done && ((spc842_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint842 = 1;
       linebuf842 = {linebuf842, spc842_phy_pc_w[8:1]};
       if (spc842_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 842, linebuf842);
          linebuf842 = "";
       end
    end else begin
       hitMadPrint842 = 0;
    end
  end
end


string linebuf843 = "";
logic hitMadPrint843 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc843_inst_done && ((spc843_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint843 = 1;
       linebuf843 = {linebuf843, spc843_phy_pc_w[8:1]};
       if (spc843_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 843, linebuf843);
          linebuf843 = "";
       end
    end else begin
       hitMadPrint843 = 0;
    end
  end
end


string linebuf844 = "";
logic hitMadPrint844 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc844_inst_done && ((spc844_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint844 = 1;
       linebuf844 = {linebuf844, spc844_phy_pc_w[8:1]};
       if (spc844_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 844, linebuf844);
          linebuf844 = "";
       end
    end else begin
       hitMadPrint844 = 0;
    end
  end
end


string linebuf845 = "";
logic hitMadPrint845 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc845_inst_done && ((spc845_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint845 = 1;
       linebuf845 = {linebuf845, spc845_phy_pc_w[8:1]};
       if (spc845_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 845, linebuf845);
          linebuf845 = "";
       end
    end else begin
       hitMadPrint845 = 0;
    end
  end
end


string linebuf846 = "";
logic hitMadPrint846 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc846_inst_done && ((spc846_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint846 = 1;
       linebuf846 = {linebuf846, spc846_phy_pc_w[8:1]};
       if (spc846_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 846, linebuf846);
          linebuf846 = "";
       end
    end else begin
       hitMadPrint846 = 0;
    end
  end
end


string linebuf847 = "";
logic hitMadPrint847 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc847_inst_done && ((spc847_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint847 = 1;
       linebuf847 = {linebuf847, spc847_phy_pc_w[8:1]};
       if (spc847_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 847, linebuf847);
          linebuf847 = "";
       end
    end else begin
       hitMadPrint847 = 0;
    end
  end
end


string linebuf848 = "";
logic hitMadPrint848 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc848_inst_done && ((spc848_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint848 = 1;
       linebuf848 = {linebuf848, spc848_phy_pc_w[8:1]};
       if (spc848_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 848, linebuf848);
          linebuf848 = "";
       end
    end else begin
       hitMadPrint848 = 0;
    end
  end
end


string linebuf849 = "";
logic hitMadPrint849 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc849_inst_done && ((spc849_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint849 = 1;
       linebuf849 = {linebuf849, spc849_phy_pc_w[8:1]};
       if (spc849_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 849, linebuf849);
          linebuf849 = "";
       end
    end else begin
       hitMadPrint849 = 0;
    end
  end
end


string linebuf850 = "";
logic hitMadPrint850 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc850_inst_done && ((spc850_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint850 = 1;
       linebuf850 = {linebuf850, spc850_phy_pc_w[8:1]};
       if (spc850_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 850, linebuf850);
          linebuf850 = "";
       end
    end else begin
       hitMadPrint850 = 0;
    end
  end
end


string linebuf851 = "";
logic hitMadPrint851 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc851_inst_done && ((spc851_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint851 = 1;
       linebuf851 = {linebuf851, spc851_phy_pc_w[8:1]};
       if (spc851_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 851, linebuf851);
          linebuf851 = "";
       end
    end else begin
       hitMadPrint851 = 0;
    end
  end
end


string linebuf852 = "";
logic hitMadPrint852 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc852_inst_done && ((spc852_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint852 = 1;
       linebuf852 = {linebuf852, spc852_phy_pc_w[8:1]};
       if (spc852_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 852, linebuf852);
          linebuf852 = "";
       end
    end else begin
       hitMadPrint852 = 0;
    end
  end
end


string linebuf853 = "";
logic hitMadPrint853 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc853_inst_done && ((spc853_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint853 = 1;
       linebuf853 = {linebuf853, spc853_phy_pc_w[8:1]};
       if (spc853_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 853, linebuf853);
          linebuf853 = "";
       end
    end else begin
       hitMadPrint853 = 0;
    end
  end
end


string linebuf854 = "";
logic hitMadPrint854 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc854_inst_done && ((spc854_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint854 = 1;
       linebuf854 = {linebuf854, spc854_phy_pc_w[8:1]};
       if (spc854_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 854, linebuf854);
          linebuf854 = "";
       end
    end else begin
       hitMadPrint854 = 0;
    end
  end
end


string linebuf855 = "";
logic hitMadPrint855 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc855_inst_done && ((spc855_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint855 = 1;
       linebuf855 = {linebuf855, spc855_phy_pc_w[8:1]};
       if (spc855_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 855, linebuf855);
          linebuf855 = "";
       end
    end else begin
       hitMadPrint855 = 0;
    end
  end
end


string linebuf856 = "";
logic hitMadPrint856 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc856_inst_done && ((spc856_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint856 = 1;
       linebuf856 = {linebuf856, spc856_phy_pc_w[8:1]};
       if (spc856_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 856, linebuf856);
          linebuf856 = "";
       end
    end else begin
       hitMadPrint856 = 0;
    end
  end
end


string linebuf857 = "";
logic hitMadPrint857 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc857_inst_done && ((spc857_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint857 = 1;
       linebuf857 = {linebuf857, spc857_phy_pc_w[8:1]};
       if (spc857_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 857, linebuf857);
          linebuf857 = "";
       end
    end else begin
       hitMadPrint857 = 0;
    end
  end
end


string linebuf858 = "";
logic hitMadPrint858 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc858_inst_done && ((spc858_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint858 = 1;
       linebuf858 = {linebuf858, spc858_phy_pc_w[8:1]};
       if (spc858_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 858, linebuf858);
          linebuf858 = "";
       end
    end else begin
       hitMadPrint858 = 0;
    end
  end
end


string linebuf859 = "";
logic hitMadPrint859 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc859_inst_done && ((spc859_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint859 = 1;
       linebuf859 = {linebuf859, spc859_phy_pc_w[8:1]};
       if (spc859_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 859, linebuf859);
          linebuf859 = "";
       end
    end else begin
       hitMadPrint859 = 0;
    end
  end
end


string linebuf860 = "";
logic hitMadPrint860 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc860_inst_done && ((spc860_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint860 = 1;
       linebuf860 = {linebuf860, spc860_phy_pc_w[8:1]};
       if (spc860_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 860, linebuf860);
          linebuf860 = "";
       end
    end else begin
       hitMadPrint860 = 0;
    end
  end
end


string linebuf861 = "";
logic hitMadPrint861 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc861_inst_done && ((spc861_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint861 = 1;
       linebuf861 = {linebuf861, spc861_phy_pc_w[8:1]};
       if (spc861_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 861, linebuf861);
          linebuf861 = "";
       end
    end else begin
       hitMadPrint861 = 0;
    end
  end
end


string linebuf862 = "";
logic hitMadPrint862 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc862_inst_done && ((spc862_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint862 = 1;
       linebuf862 = {linebuf862, spc862_phy_pc_w[8:1]};
       if (spc862_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 862, linebuf862);
          linebuf862 = "";
       end
    end else begin
       hitMadPrint862 = 0;
    end
  end
end


string linebuf863 = "";
logic hitMadPrint863 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc863_inst_done && ((spc863_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint863 = 1;
       linebuf863 = {linebuf863, spc863_phy_pc_w[8:1]};
       if (spc863_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 863, linebuf863);
          linebuf863 = "";
       end
    end else begin
       hitMadPrint863 = 0;
    end
  end
end


string linebuf864 = "";
logic hitMadPrint864 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc864_inst_done && ((spc864_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint864 = 1;
       linebuf864 = {linebuf864, spc864_phy_pc_w[8:1]};
       if (spc864_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 864, linebuf864);
          linebuf864 = "";
       end
    end else begin
       hitMadPrint864 = 0;
    end
  end
end


string linebuf865 = "";
logic hitMadPrint865 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc865_inst_done && ((spc865_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint865 = 1;
       linebuf865 = {linebuf865, spc865_phy_pc_w[8:1]};
       if (spc865_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 865, linebuf865);
          linebuf865 = "";
       end
    end else begin
       hitMadPrint865 = 0;
    end
  end
end


string linebuf866 = "";
logic hitMadPrint866 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc866_inst_done && ((spc866_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint866 = 1;
       linebuf866 = {linebuf866, spc866_phy_pc_w[8:1]};
       if (spc866_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 866, linebuf866);
          linebuf866 = "";
       end
    end else begin
       hitMadPrint866 = 0;
    end
  end
end


string linebuf867 = "";
logic hitMadPrint867 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc867_inst_done && ((spc867_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint867 = 1;
       linebuf867 = {linebuf867, spc867_phy_pc_w[8:1]};
       if (spc867_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 867, linebuf867);
          linebuf867 = "";
       end
    end else begin
       hitMadPrint867 = 0;
    end
  end
end


string linebuf868 = "";
logic hitMadPrint868 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc868_inst_done && ((spc868_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint868 = 1;
       linebuf868 = {linebuf868, spc868_phy_pc_w[8:1]};
       if (spc868_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 868, linebuf868);
          linebuf868 = "";
       end
    end else begin
       hitMadPrint868 = 0;
    end
  end
end


string linebuf869 = "";
logic hitMadPrint869 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc869_inst_done && ((spc869_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint869 = 1;
       linebuf869 = {linebuf869, spc869_phy_pc_w[8:1]};
       if (spc869_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 869, linebuf869);
          linebuf869 = "";
       end
    end else begin
       hitMadPrint869 = 0;
    end
  end
end


string linebuf870 = "";
logic hitMadPrint870 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc870_inst_done && ((spc870_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint870 = 1;
       linebuf870 = {linebuf870, spc870_phy_pc_w[8:1]};
       if (spc870_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 870, linebuf870);
          linebuf870 = "";
       end
    end else begin
       hitMadPrint870 = 0;
    end
  end
end


string linebuf871 = "";
logic hitMadPrint871 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc871_inst_done && ((spc871_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint871 = 1;
       linebuf871 = {linebuf871, spc871_phy_pc_w[8:1]};
       if (spc871_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 871, linebuf871);
          linebuf871 = "";
       end
    end else begin
       hitMadPrint871 = 0;
    end
  end
end


string linebuf872 = "";
logic hitMadPrint872 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc872_inst_done && ((spc872_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint872 = 1;
       linebuf872 = {linebuf872, spc872_phy_pc_w[8:1]};
       if (spc872_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 872, linebuf872);
          linebuf872 = "";
       end
    end else begin
       hitMadPrint872 = 0;
    end
  end
end


string linebuf873 = "";
logic hitMadPrint873 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc873_inst_done && ((spc873_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint873 = 1;
       linebuf873 = {linebuf873, spc873_phy_pc_w[8:1]};
       if (spc873_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 873, linebuf873);
          linebuf873 = "";
       end
    end else begin
       hitMadPrint873 = 0;
    end
  end
end


string linebuf874 = "";
logic hitMadPrint874 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc874_inst_done && ((spc874_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint874 = 1;
       linebuf874 = {linebuf874, spc874_phy_pc_w[8:1]};
       if (spc874_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 874, linebuf874);
          linebuf874 = "";
       end
    end else begin
       hitMadPrint874 = 0;
    end
  end
end


string linebuf875 = "";
logic hitMadPrint875 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc875_inst_done && ((spc875_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint875 = 1;
       linebuf875 = {linebuf875, spc875_phy_pc_w[8:1]};
       if (spc875_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 875, linebuf875);
          linebuf875 = "";
       end
    end else begin
       hitMadPrint875 = 0;
    end
  end
end


string linebuf876 = "";
logic hitMadPrint876 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc876_inst_done && ((spc876_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint876 = 1;
       linebuf876 = {linebuf876, spc876_phy_pc_w[8:1]};
       if (spc876_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 876, linebuf876);
          linebuf876 = "";
       end
    end else begin
       hitMadPrint876 = 0;
    end
  end
end


string linebuf877 = "";
logic hitMadPrint877 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc877_inst_done && ((spc877_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint877 = 1;
       linebuf877 = {linebuf877, spc877_phy_pc_w[8:1]};
       if (spc877_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 877, linebuf877);
          linebuf877 = "";
       end
    end else begin
       hitMadPrint877 = 0;
    end
  end
end


string linebuf878 = "";
logic hitMadPrint878 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc878_inst_done && ((spc878_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint878 = 1;
       linebuf878 = {linebuf878, spc878_phy_pc_w[8:1]};
       if (spc878_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 878, linebuf878);
          linebuf878 = "";
       end
    end else begin
       hitMadPrint878 = 0;
    end
  end
end


string linebuf879 = "";
logic hitMadPrint879 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc879_inst_done && ((spc879_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint879 = 1;
       linebuf879 = {linebuf879, spc879_phy_pc_w[8:1]};
       if (spc879_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 879, linebuf879);
          linebuf879 = "";
       end
    end else begin
       hitMadPrint879 = 0;
    end
  end
end


string linebuf880 = "";
logic hitMadPrint880 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc880_inst_done && ((spc880_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint880 = 1;
       linebuf880 = {linebuf880, spc880_phy_pc_w[8:1]};
       if (spc880_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 880, linebuf880);
          linebuf880 = "";
       end
    end else begin
       hitMadPrint880 = 0;
    end
  end
end


string linebuf881 = "";
logic hitMadPrint881 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc881_inst_done && ((spc881_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint881 = 1;
       linebuf881 = {linebuf881, spc881_phy_pc_w[8:1]};
       if (spc881_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 881, linebuf881);
          linebuf881 = "";
       end
    end else begin
       hitMadPrint881 = 0;
    end
  end
end


string linebuf882 = "";
logic hitMadPrint882 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc882_inst_done && ((spc882_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint882 = 1;
       linebuf882 = {linebuf882, spc882_phy_pc_w[8:1]};
       if (spc882_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 882, linebuf882);
          linebuf882 = "";
       end
    end else begin
       hitMadPrint882 = 0;
    end
  end
end


string linebuf883 = "";
logic hitMadPrint883 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc883_inst_done && ((spc883_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint883 = 1;
       linebuf883 = {linebuf883, spc883_phy_pc_w[8:1]};
       if (spc883_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 883, linebuf883);
          linebuf883 = "";
       end
    end else begin
       hitMadPrint883 = 0;
    end
  end
end


string linebuf884 = "";
logic hitMadPrint884 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc884_inst_done && ((spc884_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint884 = 1;
       linebuf884 = {linebuf884, spc884_phy_pc_w[8:1]};
       if (spc884_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 884, linebuf884);
          linebuf884 = "";
       end
    end else begin
       hitMadPrint884 = 0;
    end
  end
end


string linebuf885 = "";
logic hitMadPrint885 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc885_inst_done && ((spc885_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint885 = 1;
       linebuf885 = {linebuf885, spc885_phy_pc_w[8:1]};
       if (spc885_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 885, linebuf885);
          linebuf885 = "";
       end
    end else begin
       hitMadPrint885 = 0;
    end
  end
end


string linebuf886 = "";
logic hitMadPrint886 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc886_inst_done && ((spc886_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint886 = 1;
       linebuf886 = {linebuf886, spc886_phy_pc_w[8:1]};
       if (spc886_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 886, linebuf886);
          linebuf886 = "";
       end
    end else begin
       hitMadPrint886 = 0;
    end
  end
end


string linebuf887 = "";
logic hitMadPrint887 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc887_inst_done && ((spc887_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint887 = 1;
       linebuf887 = {linebuf887, spc887_phy_pc_w[8:1]};
       if (spc887_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 887, linebuf887);
          linebuf887 = "";
       end
    end else begin
       hitMadPrint887 = 0;
    end
  end
end


string linebuf888 = "";
logic hitMadPrint888 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc888_inst_done && ((spc888_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint888 = 1;
       linebuf888 = {linebuf888, spc888_phy_pc_w[8:1]};
       if (spc888_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 888, linebuf888);
          linebuf888 = "";
       end
    end else begin
       hitMadPrint888 = 0;
    end
  end
end


string linebuf889 = "";
logic hitMadPrint889 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc889_inst_done && ((spc889_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint889 = 1;
       linebuf889 = {linebuf889, spc889_phy_pc_w[8:1]};
       if (spc889_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 889, linebuf889);
          linebuf889 = "";
       end
    end else begin
       hitMadPrint889 = 0;
    end
  end
end


string linebuf890 = "";
logic hitMadPrint890 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc890_inst_done && ((spc890_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint890 = 1;
       linebuf890 = {linebuf890, spc890_phy_pc_w[8:1]};
       if (spc890_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 890, linebuf890);
          linebuf890 = "";
       end
    end else begin
       hitMadPrint890 = 0;
    end
  end
end


string linebuf891 = "";
logic hitMadPrint891 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc891_inst_done && ((spc891_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint891 = 1;
       linebuf891 = {linebuf891, spc891_phy_pc_w[8:1]};
       if (spc891_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 891, linebuf891);
          linebuf891 = "";
       end
    end else begin
       hitMadPrint891 = 0;
    end
  end
end


string linebuf892 = "";
logic hitMadPrint892 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc892_inst_done && ((spc892_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint892 = 1;
       linebuf892 = {linebuf892, spc892_phy_pc_w[8:1]};
       if (spc892_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 892, linebuf892);
          linebuf892 = "";
       end
    end else begin
       hitMadPrint892 = 0;
    end
  end
end


string linebuf893 = "";
logic hitMadPrint893 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc893_inst_done && ((spc893_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint893 = 1;
       linebuf893 = {linebuf893, spc893_phy_pc_w[8:1]};
       if (spc893_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 893, linebuf893);
          linebuf893 = "";
       end
    end else begin
       hitMadPrint893 = 0;
    end
  end
end


string linebuf894 = "";
logic hitMadPrint894 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc894_inst_done && ((spc894_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint894 = 1;
       linebuf894 = {linebuf894, spc894_phy_pc_w[8:1]};
       if (spc894_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 894, linebuf894);
          linebuf894 = "";
       end
    end else begin
       hitMadPrint894 = 0;
    end
  end
end


string linebuf895 = "";
logic hitMadPrint895 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc895_inst_done && ((spc895_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint895 = 1;
       linebuf895 = {linebuf895, spc895_phy_pc_w[8:1]};
       if (spc895_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 895, linebuf895);
          linebuf895 = "";
       end
    end else begin
       hitMadPrint895 = 0;
    end
  end
end


string linebuf896 = "";
logic hitMadPrint896 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc896_inst_done && ((spc896_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint896 = 1;
       linebuf896 = {linebuf896, spc896_phy_pc_w[8:1]};
       if (spc896_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 896, linebuf896);
          linebuf896 = "";
       end
    end else begin
       hitMadPrint896 = 0;
    end
  end
end


string linebuf897 = "";
logic hitMadPrint897 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc897_inst_done && ((spc897_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint897 = 1;
       linebuf897 = {linebuf897, spc897_phy_pc_w[8:1]};
       if (spc897_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 897, linebuf897);
          linebuf897 = "";
       end
    end else begin
       hitMadPrint897 = 0;
    end
  end
end


string linebuf898 = "";
logic hitMadPrint898 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc898_inst_done && ((spc898_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint898 = 1;
       linebuf898 = {linebuf898, spc898_phy_pc_w[8:1]};
       if (spc898_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 898, linebuf898);
          linebuf898 = "";
       end
    end else begin
       hitMadPrint898 = 0;
    end
  end
end


string linebuf899 = "";
logic hitMadPrint899 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc899_inst_done && ((spc899_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint899 = 1;
       linebuf899 = {linebuf899, spc899_phy_pc_w[8:1]};
       if (spc899_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 899, linebuf899);
          linebuf899 = "";
       end
    end else begin
       hitMadPrint899 = 0;
    end
  end
end


string linebuf900 = "";
logic hitMadPrint900 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc900_inst_done && ((spc900_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint900 = 1;
       linebuf900 = {linebuf900, spc900_phy_pc_w[8:1]};
       if (spc900_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 900, linebuf900);
          linebuf900 = "";
       end
    end else begin
       hitMadPrint900 = 0;
    end
  end
end


string linebuf901 = "";
logic hitMadPrint901 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc901_inst_done && ((spc901_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint901 = 1;
       linebuf901 = {linebuf901, spc901_phy_pc_w[8:1]};
       if (spc901_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 901, linebuf901);
          linebuf901 = "";
       end
    end else begin
       hitMadPrint901 = 0;
    end
  end
end


string linebuf902 = "";
logic hitMadPrint902 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc902_inst_done && ((spc902_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint902 = 1;
       linebuf902 = {linebuf902, spc902_phy_pc_w[8:1]};
       if (spc902_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 902, linebuf902);
          linebuf902 = "";
       end
    end else begin
       hitMadPrint902 = 0;
    end
  end
end


string linebuf903 = "";
logic hitMadPrint903 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc903_inst_done && ((spc903_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint903 = 1;
       linebuf903 = {linebuf903, spc903_phy_pc_w[8:1]};
       if (spc903_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 903, linebuf903);
          linebuf903 = "";
       end
    end else begin
       hitMadPrint903 = 0;
    end
  end
end


string linebuf904 = "";
logic hitMadPrint904 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc904_inst_done && ((spc904_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint904 = 1;
       linebuf904 = {linebuf904, spc904_phy_pc_w[8:1]};
       if (spc904_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 904, linebuf904);
          linebuf904 = "";
       end
    end else begin
       hitMadPrint904 = 0;
    end
  end
end


string linebuf905 = "";
logic hitMadPrint905 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc905_inst_done && ((spc905_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint905 = 1;
       linebuf905 = {linebuf905, spc905_phy_pc_w[8:1]};
       if (spc905_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 905, linebuf905);
          linebuf905 = "";
       end
    end else begin
       hitMadPrint905 = 0;
    end
  end
end


string linebuf906 = "";
logic hitMadPrint906 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc906_inst_done && ((spc906_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint906 = 1;
       linebuf906 = {linebuf906, spc906_phy_pc_w[8:1]};
       if (spc906_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 906, linebuf906);
          linebuf906 = "";
       end
    end else begin
       hitMadPrint906 = 0;
    end
  end
end


string linebuf907 = "";
logic hitMadPrint907 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc907_inst_done && ((spc907_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint907 = 1;
       linebuf907 = {linebuf907, spc907_phy_pc_w[8:1]};
       if (spc907_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 907, linebuf907);
          linebuf907 = "";
       end
    end else begin
       hitMadPrint907 = 0;
    end
  end
end


string linebuf908 = "";
logic hitMadPrint908 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc908_inst_done && ((spc908_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint908 = 1;
       linebuf908 = {linebuf908, spc908_phy_pc_w[8:1]};
       if (spc908_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 908, linebuf908);
          linebuf908 = "";
       end
    end else begin
       hitMadPrint908 = 0;
    end
  end
end


string linebuf909 = "";
logic hitMadPrint909 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc909_inst_done && ((spc909_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint909 = 1;
       linebuf909 = {linebuf909, spc909_phy_pc_w[8:1]};
       if (spc909_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 909, linebuf909);
          linebuf909 = "";
       end
    end else begin
       hitMadPrint909 = 0;
    end
  end
end


string linebuf910 = "";
logic hitMadPrint910 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc910_inst_done && ((spc910_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint910 = 1;
       linebuf910 = {linebuf910, spc910_phy_pc_w[8:1]};
       if (spc910_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 910, linebuf910);
          linebuf910 = "";
       end
    end else begin
       hitMadPrint910 = 0;
    end
  end
end


string linebuf911 = "";
logic hitMadPrint911 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc911_inst_done && ((spc911_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint911 = 1;
       linebuf911 = {linebuf911, spc911_phy_pc_w[8:1]};
       if (spc911_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 911, linebuf911);
          linebuf911 = "";
       end
    end else begin
       hitMadPrint911 = 0;
    end
  end
end


string linebuf912 = "";
logic hitMadPrint912 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc912_inst_done && ((spc912_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint912 = 1;
       linebuf912 = {linebuf912, spc912_phy_pc_w[8:1]};
       if (spc912_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 912, linebuf912);
          linebuf912 = "";
       end
    end else begin
       hitMadPrint912 = 0;
    end
  end
end


string linebuf913 = "";
logic hitMadPrint913 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc913_inst_done && ((spc913_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint913 = 1;
       linebuf913 = {linebuf913, spc913_phy_pc_w[8:1]};
       if (spc913_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 913, linebuf913);
          linebuf913 = "";
       end
    end else begin
       hitMadPrint913 = 0;
    end
  end
end


string linebuf914 = "";
logic hitMadPrint914 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc914_inst_done && ((spc914_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint914 = 1;
       linebuf914 = {linebuf914, spc914_phy_pc_w[8:1]};
       if (spc914_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 914, linebuf914);
          linebuf914 = "";
       end
    end else begin
       hitMadPrint914 = 0;
    end
  end
end


string linebuf915 = "";
logic hitMadPrint915 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc915_inst_done && ((spc915_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint915 = 1;
       linebuf915 = {linebuf915, spc915_phy_pc_w[8:1]};
       if (spc915_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 915, linebuf915);
          linebuf915 = "";
       end
    end else begin
       hitMadPrint915 = 0;
    end
  end
end


string linebuf916 = "";
logic hitMadPrint916 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc916_inst_done && ((spc916_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint916 = 1;
       linebuf916 = {linebuf916, spc916_phy_pc_w[8:1]};
       if (spc916_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 916, linebuf916);
          linebuf916 = "";
       end
    end else begin
       hitMadPrint916 = 0;
    end
  end
end


string linebuf917 = "";
logic hitMadPrint917 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc917_inst_done && ((spc917_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint917 = 1;
       linebuf917 = {linebuf917, spc917_phy_pc_w[8:1]};
       if (spc917_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 917, linebuf917);
          linebuf917 = "";
       end
    end else begin
       hitMadPrint917 = 0;
    end
  end
end


string linebuf918 = "";
logic hitMadPrint918 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc918_inst_done && ((spc918_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint918 = 1;
       linebuf918 = {linebuf918, spc918_phy_pc_w[8:1]};
       if (spc918_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 918, linebuf918);
          linebuf918 = "";
       end
    end else begin
       hitMadPrint918 = 0;
    end
  end
end


string linebuf919 = "";
logic hitMadPrint919 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc919_inst_done && ((spc919_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint919 = 1;
       linebuf919 = {linebuf919, spc919_phy_pc_w[8:1]};
       if (spc919_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 919, linebuf919);
          linebuf919 = "";
       end
    end else begin
       hitMadPrint919 = 0;
    end
  end
end


string linebuf920 = "";
logic hitMadPrint920 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc920_inst_done && ((spc920_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint920 = 1;
       linebuf920 = {linebuf920, spc920_phy_pc_w[8:1]};
       if (spc920_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 920, linebuf920);
          linebuf920 = "";
       end
    end else begin
       hitMadPrint920 = 0;
    end
  end
end


string linebuf921 = "";
logic hitMadPrint921 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc921_inst_done && ((spc921_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint921 = 1;
       linebuf921 = {linebuf921, spc921_phy_pc_w[8:1]};
       if (spc921_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 921, linebuf921);
          linebuf921 = "";
       end
    end else begin
       hitMadPrint921 = 0;
    end
  end
end


string linebuf922 = "";
logic hitMadPrint922 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc922_inst_done && ((spc922_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint922 = 1;
       linebuf922 = {linebuf922, spc922_phy_pc_w[8:1]};
       if (spc922_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 922, linebuf922);
          linebuf922 = "";
       end
    end else begin
       hitMadPrint922 = 0;
    end
  end
end


string linebuf923 = "";
logic hitMadPrint923 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc923_inst_done && ((spc923_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint923 = 1;
       linebuf923 = {linebuf923, spc923_phy_pc_w[8:1]};
       if (spc923_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 923, linebuf923);
          linebuf923 = "";
       end
    end else begin
       hitMadPrint923 = 0;
    end
  end
end


string linebuf924 = "";
logic hitMadPrint924 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc924_inst_done && ((spc924_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint924 = 1;
       linebuf924 = {linebuf924, spc924_phy_pc_w[8:1]};
       if (spc924_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 924, linebuf924);
          linebuf924 = "";
       end
    end else begin
       hitMadPrint924 = 0;
    end
  end
end


string linebuf925 = "";
logic hitMadPrint925 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc925_inst_done && ((spc925_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint925 = 1;
       linebuf925 = {linebuf925, spc925_phy_pc_w[8:1]};
       if (spc925_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 925, linebuf925);
          linebuf925 = "";
       end
    end else begin
       hitMadPrint925 = 0;
    end
  end
end


string linebuf926 = "";
logic hitMadPrint926 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc926_inst_done && ((spc926_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint926 = 1;
       linebuf926 = {linebuf926, spc926_phy_pc_w[8:1]};
       if (spc926_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 926, linebuf926);
          linebuf926 = "";
       end
    end else begin
       hitMadPrint926 = 0;
    end
  end
end


string linebuf927 = "";
logic hitMadPrint927 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc927_inst_done && ((spc927_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint927 = 1;
       linebuf927 = {linebuf927, spc927_phy_pc_w[8:1]};
       if (spc927_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 927, linebuf927);
          linebuf927 = "";
       end
    end else begin
       hitMadPrint927 = 0;
    end
  end
end


string linebuf928 = "";
logic hitMadPrint928 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc928_inst_done && ((spc928_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint928 = 1;
       linebuf928 = {linebuf928, spc928_phy_pc_w[8:1]};
       if (spc928_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 928, linebuf928);
          linebuf928 = "";
       end
    end else begin
       hitMadPrint928 = 0;
    end
  end
end


string linebuf929 = "";
logic hitMadPrint929 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc929_inst_done && ((spc929_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint929 = 1;
       linebuf929 = {linebuf929, spc929_phy_pc_w[8:1]};
       if (spc929_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 929, linebuf929);
          linebuf929 = "";
       end
    end else begin
       hitMadPrint929 = 0;
    end
  end
end


string linebuf930 = "";
logic hitMadPrint930 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc930_inst_done && ((spc930_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint930 = 1;
       linebuf930 = {linebuf930, spc930_phy_pc_w[8:1]};
       if (spc930_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 930, linebuf930);
          linebuf930 = "";
       end
    end else begin
       hitMadPrint930 = 0;
    end
  end
end


string linebuf931 = "";
logic hitMadPrint931 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc931_inst_done && ((spc931_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint931 = 1;
       linebuf931 = {linebuf931, spc931_phy_pc_w[8:1]};
       if (spc931_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 931, linebuf931);
          linebuf931 = "";
       end
    end else begin
       hitMadPrint931 = 0;
    end
  end
end


string linebuf932 = "";
logic hitMadPrint932 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc932_inst_done && ((spc932_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint932 = 1;
       linebuf932 = {linebuf932, spc932_phy_pc_w[8:1]};
       if (spc932_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 932, linebuf932);
          linebuf932 = "";
       end
    end else begin
       hitMadPrint932 = 0;
    end
  end
end


string linebuf933 = "";
logic hitMadPrint933 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc933_inst_done && ((spc933_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint933 = 1;
       linebuf933 = {linebuf933, spc933_phy_pc_w[8:1]};
       if (spc933_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 933, linebuf933);
          linebuf933 = "";
       end
    end else begin
       hitMadPrint933 = 0;
    end
  end
end


string linebuf934 = "";
logic hitMadPrint934 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc934_inst_done && ((spc934_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint934 = 1;
       linebuf934 = {linebuf934, spc934_phy_pc_w[8:1]};
       if (spc934_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 934, linebuf934);
          linebuf934 = "";
       end
    end else begin
       hitMadPrint934 = 0;
    end
  end
end


string linebuf935 = "";
logic hitMadPrint935 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc935_inst_done && ((spc935_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint935 = 1;
       linebuf935 = {linebuf935, spc935_phy_pc_w[8:1]};
       if (spc935_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 935, linebuf935);
          linebuf935 = "";
       end
    end else begin
       hitMadPrint935 = 0;
    end
  end
end


string linebuf936 = "";
logic hitMadPrint936 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc936_inst_done && ((spc936_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint936 = 1;
       linebuf936 = {linebuf936, spc936_phy_pc_w[8:1]};
       if (spc936_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 936, linebuf936);
          linebuf936 = "";
       end
    end else begin
       hitMadPrint936 = 0;
    end
  end
end


string linebuf937 = "";
logic hitMadPrint937 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc937_inst_done && ((spc937_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint937 = 1;
       linebuf937 = {linebuf937, spc937_phy_pc_w[8:1]};
       if (spc937_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 937, linebuf937);
          linebuf937 = "";
       end
    end else begin
       hitMadPrint937 = 0;
    end
  end
end


string linebuf938 = "";
logic hitMadPrint938 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc938_inst_done && ((spc938_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint938 = 1;
       linebuf938 = {linebuf938, spc938_phy_pc_w[8:1]};
       if (spc938_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 938, linebuf938);
          linebuf938 = "";
       end
    end else begin
       hitMadPrint938 = 0;
    end
  end
end


string linebuf939 = "";
logic hitMadPrint939 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc939_inst_done && ((spc939_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint939 = 1;
       linebuf939 = {linebuf939, spc939_phy_pc_w[8:1]};
       if (spc939_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 939, linebuf939);
          linebuf939 = "";
       end
    end else begin
       hitMadPrint939 = 0;
    end
  end
end


string linebuf940 = "";
logic hitMadPrint940 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc940_inst_done && ((spc940_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint940 = 1;
       linebuf940 = {linebuf940, spc940_phy_pc_w[8:1]};
       if (spc940_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 940, linebuf940);
          linebuf940 = "";
       end
    end else begin
       hitMadPrint940 = 0;
    end
  end
end


string linebuf941 = "";
logic hitMadPrint941 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc941_inst_done && ((spc941_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint941 = 1;
       linebuf941 = {linebuf941, spc941_phy_pc_w[8:1]};
       if (spc941_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 941, linebuf941);
          linebuf941 = "";
       end
    end else begin
       hitMadPrint941 = 0;
    end
  end
end


string linebuf942 = "";
logic hitMadPrint942 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc942_inst_done && ((spc942_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint942 = 1;
       linebuf942 = {linebuf942, spc942_phy_pc_w[8:1]};
       if (spc942_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 942, linebuf942);
          linebuf942 = "";
       end
    end else begin
       hitMadPrint942 = 0;
    end
  end
end


string linebuf943 = "";
logic hitMadPrint943 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc943_inst_done && ((spc943_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint943 = 1;
       linebuf943 = {linebuf943, spc943_phy_pc_w[8:1]};
       if (spc943_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 943, linebuf943);
          linebuf943 = "";
       end
    end else begin
       hitMadPrint943 = 0;
    end
  end
end


string linebuf944 = "";
logic hitMadPrint944 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc944_inst_done && ((spc944_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint944 = 1;
       linebuf944 = {linebuf944, spc944_phy_pc_w[8:1]};
       if (spc944_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 944, linebuf944);
          linebuf944 = "";
       end
    end else begin
       hitMadPrint944 = 0;
    end
  end
end


string linebuf945 = "";
logic hitMadPrint945 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc945_inst_done && ((spc945_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint945 = 1;
       linebuf945 = {linebuf945, spc945_phy_pc_w[8:1]};
       if (spc945_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 945, linebuf945);
          linebuf945 = "";
       end
    end else begin
       hitMadPrint945 = 0;
    end
  end
end


string linebuf946 = "";
logic hitMadPrint946 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc946_inst_done && ((spc946_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint946 = 1;
       linebuf946 = {linebuf946, spc946_phy_pc_w[8:1]};
       if (spc946_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 946, linebuf946);
          linebuf946 = "";
       end
    end else begin
       hitMadPrint946 = 0;
    end
  end
end


string linebuf947 = "";
logic hitMadPrint947 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc947_inst_done && ((spc947_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint947 = 1;
       linebuf947 = {linebuf947, spc947_phy_pc_w[8:1]};
       if (spc947_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 947, linebuf947);
          linebuf947 = "";
       end
    end else begin
       hitMadPrint947 = 0;
    end
  end
end


string linebuf948 = "";
logic hitMadPrint948 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc948_inst_done && ((spc948_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint948 = 1;
       linebuf948 = {linebuf948, spc948_phy_pc_w[8:1]};
       if (spc948_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 948, linebuf948);
          linebuf948 = "";
       end
    end else begin
       hitMadPrint948 = 0;
    end
  end
end


string linebuf949 = "";
logic hitMadPrint949 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc949_inst_done && ((spc949_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint949 = 1;
       linebuf949 = {linebuf949, spc949_phy_pc_w[8:1]};
       if (spc949_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 949, linebuf949);
          linebuf949 = "";
       end
    end else begin
       hitMadPrint949 = 0;
    end
  end
end


string linebuf950 = "";
logic hitMadPrint950 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc950_inst_done && ((spc950_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint950 = 1;
       linebuf950 = {linebuf950, spc950_phy_pc_w[8:1]};
       if (spc950_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 950, linebuf950);
          linebuf950 = "";
       end
    end else begin
       hitMadPrint950 = 0;
    end
  end
end


string linebuf951 = "";
logic hitMadPrint951 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc951_inst_done && ((spc951_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint951 = 1;
       linebuf951 = {linebuf951, spc951_phy_pc_w[8:1]};
       if (spc951_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 951, linebuf951);
          linebuf951 = "";
       end
    end else begin
       hitMadPrint951 = 0;
    end
  end
end


string linebuf952 = "";
logic hitMadPrint952 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc952_inst_done && ((spc952_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint952 = 1;
       linebuf952 = {linebuf952, spc952_phy_pc_w[8:1]};
       if (spc952_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 952, linebuf952);
          linebuf952 = "";
       end
    end else begin
       hitMadPrint952 = 0;
    end
  end
end


string linebuf953 = "";
logic hitMadPrint953 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc953_inst_done && ((spc953_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint953 = 1;
       linebuf953 = {linebuf953, spc953_phy_pc_w[8:1]};
       if (spc953_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 953, linebuf953);
          linebuf953 = "";
       end
    end else begin
       hitMadPrint953 = 0;
    end
  end
end


string linebuf954 = "";
logic hitMadPrint954 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc954_inst_done && ((spc954_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint954 = 1;
       linebuf954 = {linebuf954, spc954_phy_pc_w[8:1]};
       if (spc954_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 954, linebuf954);
          linebuf954 = "";
       end
    end else begin
       hitMadPrint954 = 0;
    end
  end
end


string linebuf955 = "";
logic hitMadPrint955 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc955_inst_done && ((spc955_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint955 = 1;
       linebuf955 = {linebuf955, spc955_phy_pc_w[8:1]};
       if (spc955_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 955, linebuf955);
          linebuf955 = "";
       end
    end else begin
       hitMadPrint955 = 0;
    end
  end
end


string linebuf956 = "";
logic hitMadPrint956 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc956_inst_done && ((spc956_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint956 = 1;
       linebuf956 = {linebuf956, spc956_phy_pc_w[8:1]};
       if (spc956_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 956, linebuf956);
          linebuf956 = "";
       end
    end else begin
       hitMadPrint956 = 0;
    end
  end
end


string linebuf957 = "";
logic hitMadPrint957 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc957_inst_done && ((spc957_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint957 = 1;
       linebuf957 = {linebuf957, spc957_phy_pc_w[8:1]};
       if (spc957_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 957, linebuf957);
          linebuf957 = "";
       end
    end else begin
       hitMadPrint957 = 0;
    end
  end
end


string linebuf958 = "";
logic hitMadPrint958 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc958_inst_done && ((spc958_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint958 = 1;
       linebuf958 = {linebuf958, spc958_phy_pc_w[8:1]};
       if (spc958_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 958, linebuf958);
          linebuf958 = "";
       end
    end else begin
       hitMadPrint958 = 0;
    end
  end
end


string linebuf959 = "";
logic hitMadPrint959 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc959_inst_done && ((spc959_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint959 = 1;
       linebuf959 = {linebuf959, spc959_phy_pc_w[8:1]};
       if (spc959_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 959, linebuf959);
          linebuf959 = "";
       end
    end else begin
       hitMadPrint959 = 0;
    end
  end
end


string linebuf960 = "";
logic hitMadPrint960 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc960_inst_done && ((spc960_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint960 = 1;
       linebuf960 = {linebuf960, spc960_phy_pc_w[8:1]};
       if (spc960_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 960, linebuf960);
          linebuf960 = "";
       end
    end else begin
       hitMadPrint960 = 0;
    end
  end
end


string linebuf961 = "";
logic hitMadPrint961 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc961_inst_done && ((spc961_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint961 = 1;
       linebuf961 = {linebuf961, spc961_phy_pc_w[8:1]};
       if (spc961_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 961, linebuf961);
          linebuf961 = "";
       end
    end else begin
       hitMadPrint961 = 0;
    end
  end
end


string linebuf962 = "";
logic hitMadPrint962 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc962_inst_done && ((spc962_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint962 = 1;
       linebuf962 = {linebuf962, spc962_phy_pc_w[8:1]};
       if (spc962_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 962, linebuf962);
          linebuf962 = "";
       end
    end else begin
       hitMadPrint962 = 0;
    end
  end
end


string linebuf963 = "";
logic hitMadPrint963 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc963_inst_done && ((spc963_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint963 = 1;
       linebuf963 = {linebuf963, spc963_phy_pc_w[8:1]};
       if (spc963_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 963, linebuf963);
          linebuf963 = "";
       end
    end else begin
       hitMadPrint963 = 0;
    end
  end
end


string linebuf964 = "";
logic hitMadPrint964 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc964_inst_done && ((spc964_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint964 = 1;
       linebuf964 = {linebuf964, spc964_phy_pc_w[8:1]};
       if (spc964_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 964, linebuf964);
          linebuf964 = "";
       end
    end else begin
       hitMadPrint964 = 0;
    end
  end
end


string linebuf965 = "";
logic hitMadPrint965 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc965_inst_done && ((spc965_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint965 = 1;
       linebuf965 = {linebuf965, spc965_phy_pc_w[8:1]};
       if (spc965_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 965, linebuf965);
          linebuf965 = "";
       end
    end else begin
       hitMadPrint965 = 0;
    end
  end
end


string linebuf966 = "";
logic hitMadPrint966 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc966_inst_done && ((spc966_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint966 = 1;
       linebuf966 = {linebuf966, spc966_phy_pc_w[8:1]};
       if (spc966_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 966, linebuf966);
          linebuf966 = "";
       end
    end else begin
       hitMadPrint966 = 0;
    end
  end
end


string linebuf967 = "";
logic hitMadPrint967 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc967_inst_done && ((spc967_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint967 = 1;
       linebuf967 = {linebuf967, spc967_phy_pc_w[8:1]};
       if (spc967_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 967, linebuf967);
          linebuf967 = "";
       end
    end else begin
       hitMadPrint967 = 0;
    end
  end
end


string linebuf968 = "";
logic hitMadPrint968 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc968_inst_done && ((spc968_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint968 = 1;
       linebuf968 = {linebuf968, spc968_phy_pc_w[8:1]};
       if (spc968_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 968, linebuf968);
          linebuf968 = "";
       end
    end else begin
       hitMadPrint968 = 0;
    end
  end
end


string linebuf969 = "";
logic hitMadPrint969 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc969_inst_done && ((spc969_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint969 = 1;
       linebuf969 = {linebuf969, spc969_phy_pc_w[8:1]};
       if (spc969_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 969, linebuf969);
          linebuf969 = "";
       end
    end else begin
       hitMadPrint969 = 0;
    end
  end
end


string linebuf970 = "";
logic hitMadPrint970 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc970_inst_done && ((spc970_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint970 = 1;
       linebuf970 = {linebuf970, spc970_phy_pc_w[8:1]};
       if (spc970_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 970, linebuf970);
          linebuf970 = "";
       end
    end else begin
       hitMadPrint970 = 0;
    end
  end
end


string linebuf971 = "";
logic hitMadPrint971 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc971_inst_done && ((spc971_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint971 = 1;
       linebuf971 = {linebuf971, spc971_phy_pc_w[8:1]};
       if (spc971_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 971, linebuf971);
          linebuf971 = "";
       end
    end else begin
       hitMadPrint971 = 0;
    end
  end
end


string linebuf972 = "";
logic hitMadPrint972 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc972_inst_done && ((spc972_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint972 = 1;
       linebuf972 = {linebuf972, spc972_phy_pc_w[8:1]};
       if (spc972_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 972, linebuf972);
          linebuf972 = "";
       end
    end else begin
       hitMadPrint972 = 0;
    end
  end
end


string linebuf973 = "";
logic hitMadPrint973 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc973_inst_done && ((spc973_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint973 = 1;
       linebuf973 = {linebuf973, spc973_phy_pc_w[8:1]};
       if (spc973_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 973, linebuf973);
          linebuf973 = "";
       end
    end else begin
       hitMadPrint973 = 0;
    end
  end
end


string linebuf974 = "";
logic hitMadPrint974 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc974_inst_done && ((spc974_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint974 = 1;
       linebuf974 = {linebuf974, spc974_phy_pc_w[8:1]};
       if (spc974_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 974, linebuf974);
          linebuf974 = "";
       end
    end else begin
       hitMadPrint974 = 0;
    end
  end
end


string linebuf975 = "";
logic hitMadPrint975 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc975_inst_done && ((spc975_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint975 = 1;
       linebuf975 = {linebuf975, spc975_phy_pc_w[8:1]};
       if (spc975_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 975, linebuf975);
          linebuf975 = "";
       end
    end else begin
       hitMadPrint975 = 0;
    end
  end
end


string linebuf976 = "";
logic hitMadPrint976 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc976_inst_done && ((spc976_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint976 = 1;
       linebuf976 = {linebuf976, spc976_phy_pc_w[8:1]};
       if (spc976_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 976, linebuf976);
          linebuf976 = "";
       end
    end else begin
       hitMadPrint976 = 0;
    end
  end
end


string linebuf977 = "";
logic hitMadPrint977 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc977_inst_done && ((spc977_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint977 = 1;
       linebuf977 = {linebuf977, spc977_phy_pc_w[8:1]};
       if (spc977_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 977, linebuf977);
          linebuf977 = "";
       end
    end else begin
       hitMadPrint977 = 0;
    end
  end
end


string linebuf978 = "";
logic hitMadPrint978 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc978_inst_done && ((spc978_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint978 = 1;
       linebuf978 = {linebuf978, spc978_phy_pc_w[8:1]};
       if (spc978_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 978, linebuf978);
          linebuf978 = "";
       end
    end else begin
       hitMadPrint978 = 0;
    end
  end
end


string linebuf979 = "";
logic hitMadPrint979 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc979_inst_done && ((spc979_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint979 = 1;
       linebuf979 = {linebuf979, spc979_phy_pc_w[8:1]};
       if (spc979_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 979, linebuf979);
          linebuf979 = "";
       end
    end else begin
       hitMadPrint979 = 0;
    end
  end
end


string linebuf980 = "";
logic hitMadPrint980 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc980_inst_done && ((spc980_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint980 = 1;
       linebuf980 = {linebuf980, spc980_phy_pc_w[8:1]};
       if (spc980_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 980, linebuf980);
          linebuf980 = "";
       end
    end else begin
       hitMadPrint980 = 0;
    end
  end
end


string linebuf981 = "";
logic hitMadPrint981 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc981_inst_done && ((spc981_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint981 = 1;
       linebuf981 = {linebuf981, spc981_phy_pc_w[8:1]};
       if (spc981_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 981, linebuf981);
          linebuf981 = "";
       end
    end else begin
       hitMadPrint981 = 0;
    end
  end
end


string linebuf982 = "";
logic hitMadPrint982 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc982_inst_done && ((spc982_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint982 = 1;
       linebuf982 = {linebuf982, spc982_phy_pc_w[8:1]};
       if (spc982_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 982, linebuf982);
          linebuf982 = "";
       end
    end else begin
       hitMadPrint982 = 0;
    end
  end
end


string linebuf983 = "";
logic hitMadPrint983 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc983_inst_done && ((spc983_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint983 = 1;
       linebuf983 = {linebuf983, spc983_phy_pc_w[8:1]};
       if (spc983_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 983, linebuf983);
          linebuf983 = "";
       end
    end else begin
       hitMadPrint983 = 0;
    end
  end
end


string linebuf984 = "";
logic hitMadPrint984 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc984_inst_done && ((spc984_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint984 = 1;
       linebuf984 = {linebuf984, spc984_phy_pc_w[8:1]};
       if (spc984_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 984, linebuf984);
          linebuf984 = "";
       end
    end else begin
       hitMadPrint984 = 0;
    end
  end
end


string linebuf985 = "";
logic hitMadPrint985 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc985_inst_done && ((spc985_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint985 = 1;
       linebuf985 = {linebuf985, spc985_phy_pc_w[8:1]};
       if (spc985_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 985, linebuf985);
          linebuf985 = "";
       end
    end else begin
       hitMadPrint985 = 0;
    end
  end
end


string linebuf986 = "";
logic hitMadPrint986 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc986_inst_done && ((spc986_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint986 = 1;
       linebuf986 = {linebuf986, spc986_phy_pc_w[8:1]};
       if (spc986_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 986, linebuf986);
          linebuf986 = "";
       end
    end else begin
       hitMadPrint986 = 0;
    end
  end
end


string linebuf987 = "";
logic hitMadPrint987 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc987_inst_done && ((spc987_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint987 = 1;
       linebuf987 = {linebuf987, spc987_phy_pc_w[8:1]};
       if (spc987_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 987, linebuf987);
          linebuf987 = "";
       end
    end else begin
       hitMadPrint987 = 0;
    end
  end
end


string linebuf988 = "";
logic hitMadPrint988 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc988_inst_done && ((spc988_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint988 = 1;
       linebuf988 = {linebuf988, spc988_phy_pc_w[8:1]};
       if (spc988_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 988, linebuf988);
          linebuf988 = "";
       end
    end else begin
       hitMadPrint988 = 0;
    end
  end
end


string linebuf989 = "";
logic hitMadPrint989 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc989_inst_done && ((spc989_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint989 = 1;
       linebuf989 = {linebuf989, spc989_phy_pc_w[8:1]};
       if (spc989_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 989, linebuf989);
          linebuf989 = "";
       end
    end else begin
       hitMadPrint989 = 0;
    end
  end
end


string linebuf990 = "";
logic hitMadPrint990 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc990_inst_done && ((spc990_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint990 = 1;
       linebuf990 = {linebuf990, spc990_phy_pc_w[8:1]};
       if (spc990_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 990, linebuf990);
          linebuf990 = "";
       end
    end else begin
       hitMadPrint990 = 0;
    end
  end
end


string linebuf991 = "";
logic hitMadPrint991 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc991_inst_done && ((spc991_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint991 = 1;
       linebuf991 = {linebuf991, spc991_phy_pc_w[8:1]};
       if (spc991_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 991, linebuf991);
          linebuf991 = "";
       end
    end else begin
       hitMadPrint991 = 0;
    end
  end
end


string linebuf992 = "";
logic hitMadPrint992 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc992_inst_done && ((spc992_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint992 = 1;
       linebuf992 = {linebuf992, spc992_phy_pc_w[8:1]};
       if (spc992_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 992, linebuf992);
          linebuf992 = "";
       end
    end else begin
       hitMadPrint992 = 0;
    end
  end
end


string linebuf993 = "";
logic hitMadPrint993 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc993_inst_done && ((spc993_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint993 = 1;
       linebuf993 = {linebuf993, spc993_phy_pc_w[8:1]};
       if (spc993_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 993, linebuf993);
          linebuf993 = "";
       end
    end else begin
       hitMadPrint993 = 0;
    end
  end
end


string linebuf994 = "";
logic hitMadPrint994 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc994_inst_done && ((spc994_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint994 = 1;
       linebuf994 = {linebuf994, spc994_phy_pc_w[8:1]};
       if (spc994_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 994, linebuf994);
          linebuf994 = "";
       end
    end else begin
       hitMadPrint994 = 0;
    end
  end
end


string linebuf995 = "";
logic hitMadPrint995 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc995_inst_done && ((spc995_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint995 = 1;
       linebuf995 = {linebuf995, spc995_phy_pc_w[8:1]};
       if (spc995_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 995, linebuf995);
          linebuf995 = "";
       end
    end else begin
       hitMadPrint995 = 0;
    end
  end
end


string linebuf996 = "";
logic hitMadPrint996 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc996_inst_done && ((spc996_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint996 = 1;
       linebuf996 = {linebuf996, spc996_phy_pc_w[8:1]};
       if (spc996_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 996, linebuf996);
          linebuf996 = "";
       end
    end else begin
       hitMadPrint996 = 0;
    end
  end
end


string linebuf997 = "";
logic hitMadPrint997 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc997_inst_done && ((spc997_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint997 = 1;
       linebuf997 = {linebuf997, spc997_phy_pc_w[8:1]};
       if (spc997_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 997, linebuf997);
          linebuf997 = "";
       end
    end else begin
       hitMadPrint997 = 0;
    end
  end
end


string linebuf998 = "";
logic hitMadPrint998 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc998_inst_done && ((spc998_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint998 = 1;
       linebuf998 = {linebuf998, spc998_phy_pc_w[8:1]};
       if (spc998_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 998, linebuf998);
          linebuf998 = "";
       end
    end else begin
       hitMadPrint998 = 0;
    end
  end
end


string linebuf999 = "";
logic hitMadPrint999 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc999_inst_done && ((spc999_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint999 = 1;
       linebuf999 = {linebuf999, spc999_phy_pc_w[8:1]};
       if (spc999_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 999, linebuf999);
          linebuf999 = "";
       end
    end else begin
       hitMadPrint999 = 0;
    end
  end
end


string linebuf1000 = "";
logic hitMadPrint1000 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc1000_inst_done && ((spc1000_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint1000 = 1;
       linebuf1000 = {linebuf1000, spc1000_phy_pc_w[8:1]};
       if (spc1000_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 1000, linebuf1000);
          linebuf1000 = "";
       end
    end else begin
       hitMadPrint1000 = 0;
    end
  end
end


string linebuf1001 = "";
logic hitMadPrint1001 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc1001_inst_done && ((spc1001_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint1001 = 1;
       linebuf1001 = {linebuf1001, spc1001_phy_pc_w[8:1]};
       if (spc1001_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 1001, linebuf1001);
          linebuf1001 = "";
       end
    end else begin
       hitMadPrint1001 = 0;
    end
  end
end


string linebuf1002 = "";
logic hitMadPrint1002 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc1002_inst_done && ((spc1002_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint1002 = 1;
       linebuf1002 = {linebuf1002, spc1002_phy_pc_w[8:1]};
       if (spc1002_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 1002, linebuf1002);
          linebuf1002 = "";
       end
    end else begin
       hitMadPrint1002 = 0;
    end
  end
end


string linebuf1003 = "";
logic hitMadPrint1003 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc1003_inst_done && ((spc1003_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint1003 = 1;
       linebuf1003 = {linebuf1003, spc1003_phy_pc_w[8:1]};
       if (spc1003_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 1003, linebuf1003);
          linebuf1003 = "";
       end
    end else begin
       hitMadPrint1003 = 0;
    end
  end
end


string linebuf1004 = "";
logic hitMadPrint1004 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc1004_inst_done && ((spc1004_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint1004 = 1;
       linebuf1004 = {linebuf1004, spc1004_phy_pc_w[8:1]};
       if (spc1004_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 1004, linebuf1004);
          linebuf1004 = "";
       end
    end else begin
       hitMadPrint1004 = 0;
    end
  end
end


string linebuf1005 = "";
logic hitMadPrint1005 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc1005_inst_done && ((spc1005_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint1005 = 1;
       linebuf1005 = {linebuf1005, spc1005_phy_pc_w[8:1]};
       if (spc1005_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 1005, linebuf1005);
          linebuf1005 = "";
       end
    end else begin
       hitMadPrint1005 = 0;
    end
  end
end


string linebuf1006 = "";
logic hitMadPrint1006 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc1006_inst_done && ((spc1006_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint1006 = 1;
       linebuf1006 = {linebuf1006, spc1006_phy_pc_w[8:1]};
       if (spc1006_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 1006, linebuf1006);
          linebuf1006 = "";
       end
    end else begin
       hitMadPrint1006 = 0;
    end
  end
end


string linebuf1007 = "";
logic hitMadPrint1007 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc1007_inst_done && ((spc1007_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint1007 = 1;
       linebuf1007 = {linebuf1007, spc1007_phy_pc_w[8:1]};
       if (spc1007_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 1007, linebuf1007);
          linebuf1007 = "";
       end
    end else begin
       hitMadPrint1007 = 0;
    end
  end
end


string linebuf1008 = "";
logic hitMadPrint1008 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc1008_inst_done && ((spc1008_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint1008 = 1;
       linebuf1008 = {linebuf1008, spc1008_phy_pc_w[8:1]};
       if (spc1008_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 1008, linebuf1008);
          linebuf1008 = "";
       end
    end else begin
       hitMadPrint1008 = 0;
    end
  end
end


string linebuf1009 = "";
logic hitMadPrint1009 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc1009_inst_done && ((spc1009_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint1009 = 1;
       linebuf1009 = {linebuf1009, spc1009_phy_pc_w[8:1]};
       if (spc1009_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 1009, linebuf1009);
          linebuf1009 = "";
       end
    end else begin
       hitMadPrint1009 = 0;
    end
  end
end


string linebuf1010 = "";
logic hitMadPrint1010 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc1010_inst_done && ((spc1010_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint1010 = 1;
       linebuf1010 = {linebuf1010, spc1010_phy_pc_w[8:1]};
       if (spc1010_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 1010, linebuf1010);
          linebuf1010 = "";
       end
    end else begin
       hitMadPrint1010 = 0;
    end
  end
end


string linebuf1011 = "";
logic hitMadPrint1011 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc1011_inst_done && ((spc1011_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint1011 = 1;
       linebuf1011 = {linebuf1011, spc1011_phy_pc_w[8:1]};
       if (spc1011_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 1011, linebuf1011);
          linebuf1011 = "";
       end
    end else begin
       hitMadPrint1011 = 0;
    end
  end
end


string linebuf1012 = "";
logic hitMadPrint1012 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc1012_inst_done && ((spc1012_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint1012 = 1;
       linebuf1012 = {linebuf1012, spc1012_phy_pc_w[8:1]};
       if (spc1012_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 1012, linebuf1012);
          linebuf1012 = "";
       end
    end else begin
       hitMadPrint1012 = 0;
    end
  end
end


string linebuf1013 = "";
logic hitMadPrint1013 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc1013_inst_done && ((spc1013_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint1013 = 1;
       linebuf1013 = {linebuf1013, spc1013_phy_pc_w[8:1]};
       if (spc1013_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 1013, linebuf1013);
          linebuf1013 = "";
       end
    end else begin
       hitMadPrint1013 = 0;
    end
  end
end


string linebuf1014 = "";
logic hitMadPrint1014 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc1014_inst_done && ((spc1014_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint1014 = 1;
       linebuf1014 = {linebuf1014, spc1014_phy_pc_w[8:1]};
       if (spc1014_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 1014, linebuf1014);
          linebuf1014 = "";
       end
    end else begin
       hitMadPrint1014 = 0;
    end
  end
end


string linebuf1015 = "";
logic hitMadPrint1015 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc1015_inst_done && ((spc1015_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint1015 = 1;
       linebuf1015 = {linebuf1015, spc1015_phy_pc_w[8:1]};
       if (spc1015_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 1015, linebuf1015);
          linebuf1015 = "";
       end
    end else begin
       hitMadPrint1015 = 0;
    end
  end
end


string linebuf1016 = "";
logic hitMadPrint1016 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc1016_inst_done && ((spc1016_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint1016 = 1;
       linebuf1016 = {linebuf1016, spc1016_phy_pc_w[8:1]};
       if (spc1016_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 1016, linebuf1016);
          linebuf1016 = "";
       end
    end else begin
       hitMadPrint1016 = 0;
    end
  end
end


string linebuf1017 = "";
logic hitMadPrint1017 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc1017_inst_done && ((spc1017_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint1017 = 1;
       linebuf1017 = {linebuf1017, spc1017_phy_pc_w[8:1]};
       if (spc1017_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 1017, linebuf1017);
          linebuf1017 = "";
       end
    end else begin
       hitMadPrint1017 = 0;
    end
  end
end


string linebuf1018 = "";
logic hitMadPrint1018 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc1018_inst_done && ((spc1018_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint1018 = 1;
       linebuf1018 = {linebuf1018, spc1018_phy_pc_w[8:1]};
       if (spc1018_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 1018, linebuf1018);
          linebuf1018 = "";
       end
    end else begin
       hitMadPrint1018 = 0;
    end
  end
end


string linebuf1019 = "";
logic hitMadPrint1019 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc1019_inst_done && ((spc1019_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint1019 = 1;
       linebuf1019 = {linebuf1019, spc1019_phy_pc_w[8:1]};
       if (spc1019_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 1019, linebuf1019);
          linebuf1019 = "";
       end
    end else begin
       hitMadPrint1019 = 0;
    end
  end
end


string linebuf1020 = "";
logic hitMadPrint1020 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc1020_inst_done && ((spc1020_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint1020 = 1;
       linebuf1020 = {linebuf1020, spc1020_phy_pc_w[8:1]};
       if (spc1020_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 1020, linebuf1020);
          linebuf1020 = "";
       end
    end else begin
       hitMadPrint1020 = 0;
    end
  end
end


string linebuf1021 = "";
logic hitMadPrint1021 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc1021_inst_done && ((spc1021_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint1021 = 1;
       linebuf1021 = {linebuf1021, spc1021_phy_pc_w[8:1]};
       if (spc1021_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 1021, linebuf1021);
          linebuf1021 = "";
       end
    end else begin
       hitMadPrint1021 = 0;
    end
  end
end


string linebuf1022 = "";
logic hitMadPrint1022 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc1022_inst_done && ((spc1022_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint1022 = 1;
       linebuf1022 = {linebuf1022, spc1022_phy_pc_w[8:1]};
       if (spc1022_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 1022, linebuf1022);
          linebuf1022 = "";
       end
    end else begin
       hitMadPrint1022 = 0;
    end
  end
end


string linebuf1023 = "";
logic hitMadPrint1023 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc1023_inst_done && ((spc1023_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint1023 = 1;
       linebuf1023 = {linebuf1023, spc1023_phy_pc_w[8:1]};
       if (spc1023_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 1023, linebuf1023);
          linebuf1023 = "";
       end
    end else begin
       hitMadPrint1023 = 0;
    end
  end
end




//main routine of pc cmp to finish the simulation.
always @(posedge clk)begin
    if(rst_l)begin
        if(|done[`PITON_NUM_TILES-1:0]) begin

        if (done[0]) begin
            timeout[long_cpuid0] = 0;
            //check_bad_trap(spc0_phy_pc_w, 0, long_cpuid0);
            if(active_thread[long_cpuid0])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc0_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid0/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 0 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid0]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc0_phy_pc_w))
                begin
                    if(good[long_cpuid0/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid0 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid0/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid0])
        end // if (done[0])

        if (done[1]) begin
            timeout[long_cpuid1] = 0;
            //check_bad_trap(spc1_phy_pc_w, 1, long_cpuid1);
            if(active_thread[long_cpuid1])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc1_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid1/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 1 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid1]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc1_phy_pc_w))
                begin
                    if(good[long_cpuid1/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid1 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid1/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid1])
        end // if (done[1])

        if (done[2]) begin
            timeout[long_cpuid2] = 0;
            //check_bad_trap(spc2_phy_pc_w, 2, long_cpuid2);
            if(active_thread[long_cpuid2])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc2_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid2/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 2 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid2]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc2_phy_pc_w))
                begin
                    if(good[long_cpuid2/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid2 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid2/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid2])
        end // if (done[2])

        if (done[3]) begin
            timeout[long_cpuid3] = 0;
            //check_bad_trap(spc3_phy_pc_w, 3, long_cpuid3);
            if(active_thread[long_cpuid3])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc3_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid3/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 3 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid3]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc3_phy_pc_w))
                begin
                    if(good[long_cpuid3/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid3 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid3/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid3])
        end // if (done[3])

        if (done[4]) begin
            timeout[long_cpuid4] = 0;
            //check_bad_trap(spc4_phy_pc_w, 4, long_cpuid4);
            if(active_thread[long_cpuid4])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc4_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid4/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 4 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid4]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc4_phy_pc_w))
                begin
                    if(good[long_cpuid4/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid4 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid4/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid4])
        end // if (done[4])

        if (done[5]) begin
            timeout[long_cpuid5] = 0;
            //check_bad_trap(spc5_phy_pc_w, 5, long_cpuid5);
            if(active_thread[long_cpuid5])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc5_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid5/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 5 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid5]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc5_phy_pc_w))
                begin
                    if(good[long_cpuid5/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid5 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid5/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid5])
        end // if (done[5])

        if (done[6]) begin
            timeout[long_cpuid6] = 0;
            //check_bad_trap(spc6_phy_pc_w, 6, long_cpuid6);
            if(active_thread[long_cpuid6])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc6_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid6/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 6 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid6]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc6_phy_pc_w))
                begin
                    if(good[long_cpuid6/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid6 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid6/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid6])
        end // if (done[6])

        if (done[7]) begin
            timeout[long_cpuid7] = 0;
            //check_bad_trap(spc7_phy_pc_w, 7, long_cpuid7);
            if(active_thread[long_cpuid7])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc7_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid7/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 7 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid7]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc7_phy_pc_w))
                begin
                    if(good[long_cpuid7/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid7 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid7/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid7])
        end // if (done[7])

        if (done[8]) begin
            timeout[long_cpuid8] = 0;
            //check_bad_trap(spc8_phy_pc_w, 8, long_cpuid8);
            if(active_thread[long_cpuid8])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc8_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid8/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 8 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid8]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc8_phy_pc_w))
                begin
                    if(good[long_cpuid8/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid8 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid8/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid8])
        end // if (done[8])

        if (done[9]) begin
            timeout[long_cpuid9] = 0;
            //check_bad_trap(spc9_phy_pc_w, 9, long_cpuid9);
            if(active_thread[long_cpuid9])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc9_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid9/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 9 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid9]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc9_phy_pc_w))
                begin
                    if(good[long_cpuid9/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid9 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid9/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid9])
        end // if (done[9])

        if (done[10]) begin
            timeout[long_cpuid10] = 0;
            //check_bad_trap(spc10_phy_pc_w, 10, long_cpuid10);
            if(active_thread[long_cpuid10])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc10_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid10/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 10 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid10]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc10_phy_pc_w))
                begin
                    if(good[long_cpuid10/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid10 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid10/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid10])
        end // if (done[10])

        if (done[11]) begin
            timeout[long_cpuid11] = 0;
            //check_bad_trap(spc11_phy_pc_w, 11, long_cpuid11);
            if(active_thread[long_cpuid11])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc11_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid11/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 11 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid11]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc11_phy_pc_w))
                begin
                    if(good[long_cpuid11/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid11 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid11/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid11])
        end // if (done[11])

        if (done[12]) begin
            timeout[long_cpuid12] = 0;
            //check_bad_trap(spc12_phy_pc_w, 12, long_cpuid12);
            if(active_thread[long_cpuid12])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc12_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid12/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 12 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid12]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc12_phy_pc_w))
                begin
                    if(good[long_cpuid12/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid12 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid12/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid12])
        end // if (done[12])

        if (done[13]) begin
            timeout[long_cpuid13] = 0;
            //check_bad_trap(spc13_phy_pc_w, 13, long_cpuid13);
            if(active_thread[long_cpuid13])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc13_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid13/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 13 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid13]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc13_phy_pc_w))
                begin
                    if(good[long_cpuid13/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid13 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid13/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid13])
        end // if (done[13])

        if (done[14]) begin
            timeout[long_cpuid14] = 0;
            //check_bad_trap(spc14_phy_pc_w, 14, long_cpuid14);
            if(active_thread[long_cpuid14])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc14_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid14/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 14 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid14]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc14_phy_pc_w))
                begin
                    if(good[long_cpuid14/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid14 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid14/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid14])
        end // if (done[14])

        if (done[15]) begin
            timeout[long_cpuid15] = 0;
            //check_bad_trap(spc15_phy_pc_w, 15, long_cpuid15);
            if(active_thread[long_cpuid15])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc15_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid15/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 15 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid15]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc15_phy_pc_w))
                begin
                    if(good[long_cpuid15/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid15 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid15/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid15])
        end // if (done[15])

        if (done[16]) begin
            timeout[long_cpuid16] = 0;
            //check_bad_trap(spc16_phy_pc_w, 16, long_cpuid16);
            if(active_thread[long_cpuid16])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc16_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid16/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 16 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid16]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc16_phy_pc_w))
                begin
                    if(good[long_cpuid16/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid16 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid16/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid16])
        end // if (done[16])

        if (done[17]) begin
            timeout[long_cpuid17] = 0;
            //check_bad_trap(spc17_phy_pc_w, 17, long_cpuid17);
            if(active_thread[long_cpuid17])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc17_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid17/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 17 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid17]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc17_phy_pc_w))
                begin
                    if(good[long_cpuid17/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid17 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid17/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid17])
        end // if (done[17])

        if (done[18]) begin
            timeout[long_cpuid18] = 0;
            //check_bad_trap(spc18_phy_pc_w, 18, long_cpuid18);
            if(active_thread[long_cpuid18])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc18_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid18/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 18 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid18]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc18_phy_pc_w))
                begin
                    if(good[long_cpuid18/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid18 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid18/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid18])
        end // if (done[18])

        if (done[19]) begin
            timeout[long_cpuid19] = 0;
            //check_bad_trap(spc19_phy_pc_w, 19, long_cpuid19);
            if(active_thread[long_cpuid19])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc19_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid19/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 19 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid19]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc19_phy_pc_w))
                begin
                    if(good[long_cpuid19/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid19 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid19/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid19])
        end // if (done[19])

        if (done[20]) begin
            timeout[long_cpuid20] = 0;
            //check_bad_trap(spc20_phy_pc_w, 20, long_cpuid20);
            if(active_thread[long_cpuid20])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc20_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid20/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 20 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid20]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc20_phy_pc_w))
                begin
                    if(good[long_cpuid20/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid20 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid20/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid20])
        end // if (done[20])

        if (done[21]) begin
            timeout[long_cpuid21] = 0;
            //check_bad_trap(spc21_phy_pc_w, 21, long_cpuid21);
            if(active_thread[long_cpuid21])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc21_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid21/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 21 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid21]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc21_phy_pc_w))
                begin
                    if(good[long_cpuid21/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid21 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid21/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid21])
        end // if (done[21])

        if (done[22]) begin
            timeout[long_cpuid22] = 0;
            //check_bad_trap(spc22_phy_pc_w, 22, long_cpuid22);
            if(active_thread[long_cpuid22])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc22_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid22/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 22 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid22]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc22_phy_pc_w))
                begin
                    if(good[long_cpuid22/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid22 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid22/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid22])
        end // if (done[22])

        if (done[23]) begin
            timeout[long_cpuid23] = 0;
            //check_bad_trap(spc23_phy_pc_w, 23, long_cpuid23);
            if(active_thread[long_cpuid23])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc23_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid23/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 23 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid23]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc23_phy_pc_w))
                begin
                    if(good[long_cpuid23/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid23 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid23/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid23])
        end // if (done[23])

        if (done[24]) begin
            timeout[long_cpuid24] = 0;
            //check_bad_trap(spc24_phy_pc_w, 24, long_cpuid24);
            if(active_thread[long_cpuid24])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc24_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid24/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 24 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid24]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc24_phy_pc_w))
                begin
                    if(good[long_cpuid24/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid24 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid24/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid24])
        end // if (done[24])

        if (done[25]) begin
            timeout[long_cpuid25] = 0;
            //check_bad_trap(spc25_phy_pc_w, 25, long_cpuid25);
            if(active_thread[long_cpuid25])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc25_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid25/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 25 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid25]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc25_phy_pc_w))
                begin
                    if(good[long_cpuid25/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid25 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid25/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid25])
        end // if (done[25])

        if (done[26]) begin
            timeout[long_cpuid26] = 0;
            //check_bad_trap(spc26_phy_pc_w, 26, long_cpuid26);
            if(active_thread[long_cpuid26])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc26_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid26/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 26 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid26]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc26_phy_pc_w))
                begin
                    if(good[long_cpuid26/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid26 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid26/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid26])
        end // if (done[26])

        if (done[27]) begin
            timeout[long_cpuid27] = 0;
            //check_bad_trap(spc27_phy_pc_w, 27, long_cpuid27);
            if(active_thread[long_cpuid27])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc27_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid27/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 27 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid27]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc27_phy_pc_w))
                begin
                    if(good[long_cpuid27/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid27 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid27/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid27])
        end // if (done[27])

        if (done[28]) begin
            timeout[long_cpuid28] = 0;
            //check_bad_trap(spc28_phy_pc_w, 28, long_cpuid28);
            if(active_thread[long_cpuid28])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc28_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid28/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 28 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid28]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc28_phy_pc_w))
                begin
                    if(good[long_cpuid28/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid28 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid28/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid28])
        end // if (done[28])

        if (done[29]) begin
            timeout[long_cpuid29] = 0;
            //check_bad_trap(spc29_phy_pc_w, 29, long_cpuid29);
            if(active_thread[long_cpuid29])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc29_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid29/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 29 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid29]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc29_phy_pc_w))
                begin
                    if(good[long_cpuid29/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid29 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid29/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid29])
        end // if (done[29])

        if (done[30]) begin
            timeout[long_cpuid30] = 0;
            //check_bad_trap(spc30_phy_pc_w, 30, long_cpuid30);
            if(active_thread[long_cpuid30])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc30_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid30/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 30 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid30]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc30_phy_pc_w))
                begin
                    if(good[long_cpuid30/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid30 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid30/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid30])
        end // if (done[30])

        if (done[31]) begin
            timeout[long_cpuid31] = 0;
            //check_bad_trap(spc31_phy_pc_w, 31, long_cpuid31);
            if(active_thread[long_cpuid31])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc31_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid31/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 31 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid31]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc31_phy_pc_w))
                begin
                    if(good[long_cpuid31/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid31 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid31/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid31])
        end // if (done[31])

        if (done[32]) begin
            timeout[long_cpuid32] = 0;
            //check_bad_trap(spc32_phy_pc_w, 32, long_cpuid32);
            if(active_thread[long_cpuid32])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc32_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid32/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 32 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid32]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc32_phy_pc_w))
                begin
                    if(good[long_cpuid32/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid32 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid32/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid32])
        end // if (done[32])

        if (done[33]) begin
            timeout[long_cpuid33] = 0;
            //check_bad_trap(spc33_phy_pc_w, 33, long_cpuid33);
            if(active_thread[long_cpuid33])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc33_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid33/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 33 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid33]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc33_phy_pc_w))
                begin
                    if(good[long_cpuid33/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid33 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid33/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid33])
        end // if (done[33])

        if (done[34]) begin
            timeout[long_cpuid34] = 0;
            //check_bad_trap(spc34_phy_pc_w, 34, long_cpuid34);
            if(active_thread[long_cpuid34])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc34_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid34/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 34 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid34]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc34_phy_pc_w))
                begin
                    if(good[long_cpuid34/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid34 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid34/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid34])
        end // if (done[34])

        if (done[35]) begin
            timeout[long_cpuid35] = 0;
            //check_bad_trap(spc35_phy_pc_w, 35, long_cpuid35);
            if(active_thread[long_cpuid35])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc35_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid35/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 35 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid35]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc35_phy_pc_w))
                begin
                    if(good[long_cpuid35/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid35 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid35/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid35])
        end // if (done[35])

        if (done[36]) begin
            timeout[long_cpuid36] = 0;
            //check_bad_trap(spc36_phy_pc_w, 36, long_cpuid36);
            if(active_thread[long_cpuid36])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc36_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid36/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 36 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid36]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc36_phy_pc_w))
                begin
                    if(good[long_cpuid36/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid36 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid36/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid36])
        end // if (done[36])

        if (done[37]) begin
            timeout[long_cpuid37] = 0;
            //check_bad_trap(spc37_phy_pc_w, 37, long_cpuid37);
            if(active_thread[long_cpuid37])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc37_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid37/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 37 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid37]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc37_phy_pc_w))
                begin
                    if(good[long_cpuid37/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid37 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid37/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid37])
        end // if (done[37])

        if (done[38]) begin
            timeout[long_cpuid38] = 0;
            //check_bad_trap(spc38_phy_pc_w, 38, long_cpuid38);
            if(active_thread[long_cpuid38])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc38_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid38/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 38 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid38]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc38_phy_pc_w))
                begin
                    if(good[long_cpuid38/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid38 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid38/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid38])
        end // if (done[38])

        if (done[39]) begin
            timeout[long_cpuid39] = 0;
            //check_bad_trap(spc39_phy_pc_w, 39, long_cpuid39);
            if(active_thread[long_cpuid39])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc39_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid39/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 39 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid39]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc39_phy_pc_w))
                begin
                    if(good[long_cpuid39/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid39 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid39/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid39])
        end // if (done[39])

        if (done[40]) begin
            timeout[long_cpuid40] = 0;
            //check_bad_trap(spc40_phy_pc_w, 40, long_cpuid40);
            if(active_thread[long_cpuid40])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc40_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid40/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 40 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid40]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc40_phy_pc_w))
                begin
                    if(good[long_cpuid40/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid40 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid40/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid40])
        end // if (done[40])

        if (done[41]) begin
            timeout[long_cpuid41] = 0;
            //check_bad_trap(spc41_phy_pc_w, 41, long_cpuid41);
            if(active_thread[long_cpuid41])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc41_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid41/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 41 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid41]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc41_phy_pc_w))
                begin
                    if(good[long_cpuid41/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid41 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid41/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid41])
        end // if (done[41])

        if (done[42]) begin
            timeout[long_cpuid42] = 0;
            //check_bad_trap(spc42_phy_pc_w, 42, long_cpuid42);
            if(active_thread[long_cpuid42])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc42_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid42/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 42 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid42]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc42_phy_pc_w))
                begin
                    if(good[long_cpuid42/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid42 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid42/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid42])
        end // if (done[42])

        if (done[43]) begin
            timeout[long_cpuid43] = 0;
            //check_bad_trap(spc43_phy_pc_w, 43, long_cpuid43);
            if(active_thread[long_cpuid43])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc43_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid43/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 43 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid43]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc43_phy_pc_w))
                begin
                    if(good[long_cpuid43/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid43 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid43/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid43])
        end // if (done[43])

        if (done[44]) begin
            timeout[long_cpuid44] = 0;
            //check_bad_trap(spc44_phy_pc_w, 44, long_cpuid44);
            if(active_thread[long_cpuid44])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc44_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid44/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 44 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid44]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc44_phy_pc_w))
                begin
                    if(good[long_cpuid44/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid44 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid44/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid44])
        end // if (done[44])

        if (done[45]) begin
            timeout[long_cpuid45] = 0;
            //check_bad_trap(spc45_phy_pc_w, 45, long_cpuid45);
            if(active_thread[long_cpuid45])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc45_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid45/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 45 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid45]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc45_phy_pc_w))
                begin
                    if(good[long_cpuid45/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid45 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid45/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid45])
        end // if (done[45])

        if (done[46]) begin
            timeout[long_cpuid46] = 0;
            //check_bad_trap(spc46_phy_pc_w, 46, long_cpuid46);
            if(active_thread[long_cpuid46])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc46_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid46/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 46 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid46]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc46_phy_pc_w))
                begin
                    if(good[long_cpuid46/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid46 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid46/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid46])
        end // if (done[46])

        if (done[47]) begin
            timeout[long_cpuid47] = 0;
            //check_bad_trap(spc47_phy_pc_w, 47, long_cpuid47);
            if(active_thread[long_cpuid47])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc47_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid47/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 47 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid47]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc47_phy_pc_w))
                begin
                    if(good[long_cpuid47/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid47 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid47/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid47])
        end // if (done[47])

        if (done[48]) begin
            timeout[long_cpuid48] = 0;
            //check_bad_trap(spc48_phy_pc_w, 48, long_cpuid48);
            if(active_thread[long_cpuid48])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc48_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid48/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 48 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid48]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc48_phy_pc_w))
                begin
                    if(good[long_cpuid48/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid48 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid48/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid48])
        end // if (done[48])

        if (done[49]) begin
            timeout[long_cpuid49] = 0;
            //check_bad_trap(spc49_phy_pc_w, 49, long_cpuid49);
            if(active_thread[long_cpuid49])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc49_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid49/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 49 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid49]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc49_phy_pc_w))
                begin
                    if(good[long_cpuid49/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid49 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid49/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid49])
        end // if (done[49])

        if (done[50]) begin
            timeout[long_cpuid50] = 0;
            //check_bad_trap(spc50_phy_pc_w, 50, long_cpuid50);
            if(active_thread[long_cpuid50])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc50_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid50/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 50 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid50]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc50_phy_pc_w))
                begin
                    if(good[long_cpuid50/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid50 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid50/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid50])
        end // if (done[50])

        if (done[51]) begin
            timeout[long_cpuid51] = 0;
            //check_bad_trap(spc51_phy_pc_w, 51, long_cpuid51);
            if(active_thread[long_cpuid51])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc51_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid51/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 51 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid51]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc51_phy_pc_w))
                begin
                    if(good[long_cpuid51/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid51 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid51/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid51])
        end // if (done[51])

        if (done[52]) begin
            timeout[long_cpuid52] = 0;
            //check_bad_trap(spc52_phy_pc_w, 52, long_cpuid52);
            if(active_thread[long_cpuid52])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc52_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid52/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 52 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid52]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc52_phy_pc_w))
                begin
                    if(good[long_cpuid52/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid52 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid52/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid52])
        end // if (done[52])

        if (done[53]) begin
            timeout[long_cpuid53] = 0;
            //check_bad_trap(spc53_phy_pc_w, 53, long_cpuid53);
            if(active_thread[long_cpuid53])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc53_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid53/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 53 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid53]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc53_phy_pc_w))
                begin
                    if(good[long_cpuid53/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid53 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid53/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid53])
        end // if (done[53])

        if (done[54]) begin
            timeout[long_cpuid54] = 0;
            //check_bad_trap(spc54_phy_pc_w, 54, long_cpuid54);
            if(active_thread[long_cpuid54])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc54_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid54/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 54 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid54]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc54_phy_pc_w))
                begin
                    if(good[long_cpuid54/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid54 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid54/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid54])
        end // if (done[54])

        if (done[55]) begin
            timeout[long_cpuid55] = 0;
            //check_bad_trap(spc55_phy_pc_w, 55, long_cpuid55);
            if(active_thread[long_cpuid55])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc55_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid55/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 55 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid55]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc55_phy_pc_w))
                begin
                    if(good[long_cpuid55/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid55 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid55/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid55])
        end // if (done[55])

        if (done[56]) begin
            timeout[long_cpuid56] = 0;
            //check_bad_trap(spc56_phy_pc_w, 56, long_cpuid56);
            if(active_thread[long_cpuid56])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc56_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid56/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 56 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid56]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc56_phy_pc_w))
                begin
                    if(good[long_cpuid56/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid56 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid56/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid56])
        end // if (done[56])

        if (done[57]) begin
            timeout[long_cpuid57] = 0;
            //check_bad_trap(spc57_phy_pc_w, 57, long_cpuid57);
            if(active_thread[long_cpuid57])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc57_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid57/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 57 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid57]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc57_phy_pc_w))
                begin
                    if(good[long_cpuid57/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid57 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid57/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid57])
        end // if (done[57])

        if (done[58]) begin
            timeout[long_cpuid58] = 0;
            //check_bad_trap(spc58_phy_pc_w, 58, long_cpuid58);
            if(active_thread[long_cpuid58])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc58_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid58/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 58 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid58]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc58_phy_pc_w))
                begin
                    if(good[long_cpuid58/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid58 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid58/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid58])
        end // if (done[58])

        if (done[59]) begin
            timeout[long_cpuid59] = 0;
            //check_bad_trap(spc59_phy_pc_w, 59, long_cpuid59);
            if(active_thread[long_cpuid59])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc59_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid59/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 59 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid59]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc59_phy_pc_w))
                begin
                    if(good[long_cpuid59/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid59 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid59/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid59])
        end // if (done[59])

        if (done[60]) begin
            timeout[long_cpuid60] = 0;
            //check_bad_trap(spc60_phy_pc_w, 60, long_cpuid60);
            if(active_thread[long_cpuid60])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc60_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid60/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 60 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid60]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc60_phy_pc_w))
                begin
                    if(good[long_cpuid60/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid60 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid60/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid60])
        end // if (done[60])

        if (done[61]) begin
            timeout[long_cpuid61] = 0;
            //check_bad_trap(spc61_phy_pc_w, 61, long_cpuid61);
            if(active_thread[long_cpuid61])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc61_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid61/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 61 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid61]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc61_phy_pc_w))
                begin
                    if(good[long_cpuid61/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid61 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid61/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid61])
        end // if (done[61])

        if (done[62]) begin
            timeout[long_cpuid62] = 0;
            //check_bad_trap(spc62_phy_pc_w, 62, long_cpuid62);
            if(active_thread[long_cpuid62])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc62_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid62/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 62 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid62]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc62_phy_pc_w))
                begin
                    if(good[long_cpuid62/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid62 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid62/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid62])
        end // if (done[62])

        if (done[63]) begin
            timeout[long_cpuid63] = 0;
            //check_bad_trap(spc63_phy_pc_w, 63, long_cpuid63);
            if(active_thread[long_cpuid63])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc63_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid63/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 63 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid63]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc63_phy_pc_w))
                begin
                    if(good[long_cpuid63/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid63 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid63/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid63])
        end // if (done[63])

        if (done[64]) begin
            timeout[long_cpuid64] = 0;
            //check_bad_trap(spc64_phy_pc_w, 64, long_cpuid64);
            if(active_thread[long_cpuid64])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc64_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid64/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 64 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid64]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc64_phy_pc_w))
                begin
                    if(good[long_cpuid64/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid64 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid64/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid64])
        end // if (done[64])

        if (done[65]) begin
            timeout[long_cpuid65] = 0;
            //check_bad_trap(spc65_phy_pc_w, 65, long_cpuid65);
            if(active_thread[long_cpuid65])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc65_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid65/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 65 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid65]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc65_phy_pc_w))
                begin
                    if(good[long_cpuid65/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid65 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid65/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid65])
        end // if (done[65])

        if (done[66]) begin
            timeout[long_cpuid66] = 0;
            //check_bad_trap(spc66_phy_pc_w, 66, long_cpuid66);
            if(active_thread[long_cpuid66])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc66_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid66/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 66 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid66]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc66_phy_pc_w))
                begin
                    if(good[long_cpuid66/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid66 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid66/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid66])
        end // if (done[66])

        if (done[67]) begin
            timeout[long_cpuid67] = 0;
            //check_bad_trap(spc67_phy_pc_w, 67, long_cpuid67);
            if(active_thread[long_cpuid67])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc67_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid67/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 67 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid67]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc67_phy_pc_w))
                begin
                    if(good[long_cpuid67/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid67 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid67/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid67])
        end // if (done[67])

        if (done[68]) begin
            timeout[long_cpuid68] = 0;
            //check_bad_trap(spc68_phy_pc_w, 68, long_cpuid68);
            if(active_thread[long_cpuid68])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc68_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid68/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 68 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid68]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc68_phy_pc_w))
                begin
                    if(good[long_cpuid68/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid68 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid68/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid68])
        end // if (done[68])

        if (done[69]) begin
            timeout[long_cpuid69] = 0;
            //check_bad_trap(spc69_phy_pc_w, 69, long_cpuid69);
            if(active_thread[long_cpuid69])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc69_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid69/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 69 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid69]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc69_phy_pc_w))
                begin
                    if(good[long_cpuid69/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid69 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid69/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid69])
        end // if (done[69])

        if (done[70]) begin
            timeout[long_cpuid70] = 0;
            //check_bad_trap(spc70_phy_pc_w, 70, long_cpuid70);
            if(active_thread[long_cpuid70])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc70_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid70/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 70 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid70]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc70_phy_pc_w))
                begin
                    if(good[long_cpuid70/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid70 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid70/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid70])
        end // if (done[70])

        if (done[71]) begin
            timeout[long_cpuid71] = 0;
            //check_bad_trap(spc71_phy_pc_w, 71, long_cpuid71);
            if(active_thread[long_cpuid71])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc71_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid71/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 71 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid71]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc71_phy_pc_w))
                begin
                    if(good[long_cpuid71/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid71 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid71/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid71])
        end // if (done[71])

        if (done[72]) begin
            timeout[long_cpuid72] = 0;
            //check_bad_trap(spc72_phy_pc_w, 72, long_cpuid72);
            if(active_thread[long_cpuid72])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc72_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid72/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 72 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid72]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc72_phy_pc_w))
                begin
                    if(good[long_cpuid72/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid72 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid72/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid72])
        end // if (done[72])

        if (done[73]) begin
            timeout[long_cpuid73] = 0;
            //check_bad_trap(spc73_phy_pc_w, 73, long_cpuid73);
            if(active_thread[long_cpuid73])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc73_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid73/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 73 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid73]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc73_phy_pc_w))
                begin
                    if(good[long_cpuid73/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid73 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid73/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid73])
        end // if (done[73])

        if (done[74]) begin
            timeout[long_cpuid74] = 0;
            //check_bad_trap(spc74_phy_pc_w, 74, long_cpuid74);
            if(active_thread[long_cpuid74])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc74_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid74/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 74 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid74]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc74_phy_pc_w))
                begin
                    if(good[long_cpuid74/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid74 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid74/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid74])
        end // if (done[74])

        if (done[75]) begin
            timeout[long_cpuid75] = 0;
            //check_bad_trap(spc75_phy_pc_w, 75, long_cpuid75);
            if(active_thread[long_cpuid75])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc75_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid75/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 75 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid75]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc75_phy_pc_w))
                begin
                    if(good[long_cpuid75/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid75 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid75/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid75])
        end // if (done[75])

        if (done[76]) begin
            timeout[long_cpuid76] = 0;
            //check_bad_trap(spc76_phy_pc_w, 76, long_cpuid76);
            if(active_thread[long_cpuid76])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc76_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid76/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 76 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid76]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc76_phy_pc_w))
                begin
                    if(good[long_cpuid76/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid76 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid76/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid76])
        end // if (done[76])

        if (done[77]) begin
            timeout[long_cpuid77] = 0;
            //check_bad_trap(spc77_phy_pc_w, 77, long_cpuid77);
            if(active_thread[long_cpuid77])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc77_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid77/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 77 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid77]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc77_phy_pc_w))
                begin
                    if(good[long_cpuid77/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid77 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid77/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid77])
        end // if (done[77])

        if (done[78]) begin
            timeout[long_cpuid78] = 0;
            //check_bad_trap(spc78_phy_pc_w, 78, long_cpuid78);
            if(active_thread[long_cpuid78])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc78_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid78/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 78 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid78]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc78_phy_pc_w))
                begin
                    if(good[long_cpuid78/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid78 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid78/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid78])
        end // if (done[78])

        if (done[79]) begin
            timeout[long_cpuid79] = 0;
            //check_bad_trap(spc79_phy_pc_w, 79, long_cpuid79);
            if(active_thread[long_cpuid79])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc79_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid79/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 79 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid79]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc79_phy_pc_w))
                begin
                    if(good[long_cpuid79/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid79 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid79/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid79])
        end // if (done[79])

        if (done[80]) begin
            timeout[long_cpuid80] = 0;
            //check_bad_trap(spc80_phy_pc_w, 80, long_cpuid80);
            if(active_thread[long_cpuid80])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc80_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid80/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 80 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid80]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc80_phy_pc_w))
                begin
                    if(good[long_cpuid80/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid80 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid80/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid80])
        end // if (done[80])

        if (done[81]) begin
            timeout[long_cpuid81] = 0;
            //check_bad_trap(spc81_phy_pc_w, 81, long_cpuid81);
            if(active_thread[long_cpuid81])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc81_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid81/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 81 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid81]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc81_phy_pc_w))
                begin
                    if(good[long_cpuid81/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid81 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid81/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid81])
        end // if (done[81])

        if (done[82]) begin
            timeout[long_cpuid82] = 0;
            //check_bad_trap(spc82_phy_pc_w, 82, long_cpuid82);
            if(active_thread[long_cpuid82])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc82_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid82/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 82 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid82]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc82_phy_pc_w))
                begin
                    if(good[long_cpuid82/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid82 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid82/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid82])
        end // if (done[82])

        if (done[83]) begin
            timeout[long_cpuid83] = 0;
            //check_bad_trap(spc83_phy_pc_w, 83, long_cpuid83);
            if(active_thread[long_cpuid83])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc83_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid83/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 83 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid83]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc83_phy_pc_w))
                begin
                    if(good[long_cpuid83/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid83 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid83/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid83])
        end // if (done[83])

        if (done[84]) begin
            timeout[long_cpuid84] = 0;
            //check_bad_trap(spc84_phy_pc_w, 84, long_cpuid84);
            if(active_thread[long_cpuid84])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc84_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid84/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 84 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid84]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc84_phy_pc_w))
                begin
                    if(good[long_cpuid84/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid84 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid84/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid84])
        end // if (done[84])

        if (done[85]) begin
            timeout[long_cpuid85] = 0;
            //check_bad_trap(spc85_phy_pc_w, 85, long_cpuid85);
            if(active_thread[long_cpuid85])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc85_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid85/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 85 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid85]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc85_phy_pc_w))
                begin
                    if(good[long_cpuid85/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid85 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid85/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid85])
        end // if (done[85])

        if (done[86]) begin
            timeout[long_cpuid86] = 0;
            //check_bad_trap(spc86_phy_pc_w, 86, long_cpuid86);
            if(active_thread[long_cpuid86])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc86_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid86/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 86 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid86]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc86_phy_pc_w))
                begin
                    if(good[long_cpuid86/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid86 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid86/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid86])
        end // if (done[86])

        if (done[87]) begin
            timeout[long_cpuid87] = 0;
            //check_bad_trap(spc87_phy_pc_w, 87, long_cpuid87);
            if(active_thread[long_cpuid87])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc87_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid87/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 87 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid87]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc87_phy_pc_w))
                begin
                    if(good[long_cpuid87/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid87 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid87/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid87])
        end // if (done[87])

        if (done[88]) begin
            timeout[long_cpuid88] = 0;
            //check_bad_trap(spc88_phy_pc_w, 88, long_cpuid88);
            if(active_thread[long_cpuid88])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc88_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid88/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 88 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid88]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc88_phy_pc_w))
                begin
                    if(good[long_cpuid88/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid88 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid88/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid88])
        end // if (done[88])

        if (done[89]) begin
            timeout[long_cpuid89] = 0;
            //check_bad_trap(spc89_phy_pc_w, 89, long_cpuid89);
            if(active_thread[long_cpuid89])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc89_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid89/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 89 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid89]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc89_phy_pc_w))
                begin
                    if(good[long_cpuid89/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid89 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid89/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid89])
        end // if (done[89])

        if (done[90]) begin
            timeout[long_cpuid90] = 0;
            //check_bad_trap(spc90_phy_pc_w, 90, long_cpuid90);
            if(active_thread[long_cpuid90])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc90_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid90/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 90 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid90]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc90_phy_pc_w))
                begin
                    if(good[long_cpuid90/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid90 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid90/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid90])
        end // if (done[90])

        if (done[91]) begin
            timeout[long_cpuid91] = 0;
            //check_bad_trap(spc91_phy_pc_w, 91, long_cpuid91);
            if(active_thread[long_cpuid91])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc91_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid91/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 91 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid91]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc91_phy_pc_w))
                begin
                    if(good[long_cpuid91/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid91 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid91/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid91])
        end // if (done[91])

        if (done[92]) begin
            timeout[long_cpuid92] = 0;
            //check_bad_trap(spc92_phy_pc_w, 92, long_cpuid92);
            if(active_thread[long_cpuid92])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc92_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid92/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 92 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid92]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc92_phy_pc_w))
                begin
                    if(good[long_cpuid92/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid92 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid92/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid92])
        end // if (done[92])

        if (done[93]) begin
            timeout[long_cpuid93] = 0;
            //check_bad_trap(spc93_phy_pc_w, 93, long_cpuid93);
            if(active_thread[long_cpuid93])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc93_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid93/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 93 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid93]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc93_phy_pc_w))
                begin
                    if(good[long_cpuid93/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid93 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid93/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid93])
        end // if (done[93])

        if (done[94]) begin
            timeout[long_cpuid94] = 0;
            //check_bad_trap(spc94_phy_pc_w, 94, long_cpuid94);
            if(active_thread[long_cpuid94])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc94_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid94/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 94 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid94]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc94_phy_pc_w))
                begin
                    if(good[long_cpuid94/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid94 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid94/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid94])
        end // if (done[94])

        if (done[95]) begin
            timeout[long_cpuid95] = 0;
            //check_bad_trap(spc95_phy_pc_w, 95, long_cpuid95);
            if(active_thread[long_cpuid95])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc95_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid95/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 95 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid95]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc95_phy_pc_w))
                begin
                    if(good[long_cpuid95/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid95 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid95/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid95])
        end // if (done[95])

        if (done[96]) begin
            timeout[long_cpuid96] = 0;
            //check_bad_trap(spc96_phy_pc_w, 96, long_cpuid96);
            if(active_thread[long_cpuid96])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc96_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid96/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 96 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid96]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc96_phy_pc_w))
                begin
                    if(good[long_cpuid96/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid96 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid96/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid96])
        end // if (done[96])

        if (done[97]) begin
            timeout[long_cpuid97] = 0;
            //check_bad_trap(spc97_phy_pc_w, 97, long_cpuid97);
            if(active_thread[long_cpuid97])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc97_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid97/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 97 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid97]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc97_phy_pc_w))
                begin
                    if(good[long_cpuid97/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid97 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid97/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid97])
        end // if (done[97])

        if (done[98]) begin
            timeout[long_cpuid98] = 0;
            //check_bad_trap(spc98_phy_pc_w, 98, long_cpuid98);
            if(active_thread[long_cpuid98])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc98_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid98/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 98 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid98]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc98_phy_pc_w))
                begin
                    if(good[long_cpuid98/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid98 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid98/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid98])
        end // if (done[98])

        if (done[99]) begin
            timeout[long_cpuid99] = 0;
            //check_bad_trap(spc99_phy_pc_w, 99, long_cpuid99);
            if(active_thread[long_cpuid99])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc99_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid99/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 99 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid99]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc99_phy_pc_w))
                begin
                    if(good[long_cpuid99/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid99 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid99/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid99])
        end // if (done[99])

        if (done[100]) begin
            timeout[long_cpuid100] = 0;
            //check_bad_trap(spc100_phy_pc_w, 100, long_cpuid100);
            if(active_thread[long_cpuid100])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc100_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid100/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 100 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid100]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc100_phy_pc_w))
                begin
                    if(good[long_cpuid100/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid100 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid100/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid100])
        end // if (done[100])

        if (done[101]) begin
            timeout[long_cpuid101] = 0;
            //check_bad_trap(spc101_phy_pc_w, 101, long_cpuid101);
            if(active_thread[long_cpuid101])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc101_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid101/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 101 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid101]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc101_phy_pc_w))
                begin
                    if(good[long_cpuid101/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid101 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid101/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid101])
        end // if (done[101])

        if (done[102]) begin
            timeout[long_cpuid102] = 0;
            //check_bad_trap(spc102_phy_pc_w, 102, long_cpuid102);
            if(active_thread[long_cpuid102])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc102_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid102/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 102 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid102]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc102_phy_pc_w))
                begin
                    if(good[long_cpuid102/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid102 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid102/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid102])
        end // if (done[102])

        if (done[103]) begin
            timeout[long_cpuid103] = 0;
            //check_bad_trap(spc103_phy_pc_w, 103, long_cpuid103);
            if(active_thread[long_cpuid103])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc103_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid103/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 103 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid103]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc103_phy_pc_w))
                begin
                    if(good[long_cpuid103/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid103 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid103/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid103])
        end // if (done[103])

        if (done[104]) begin
            timeout[long_cpuid104] = 0;
            //check_bad_trap(spc104_phy_pc_w, 104, long_cpuid104);
            if(active_thread[long_cpuid104])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc104_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid104/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 104 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid104]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc104_phy_pc_w))
                begin
                    if(good[long_cpuid104/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid104 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid104/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid104])
        end // if (done[104])

        if (done[105]) begin
            timeout[long_cpuid105] = 0;
            //check_bad_trap(spc105_phy_pc_w, 105, long_cpuid105);
            if(active_thread[long_cpuid105])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc105_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid105/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 105 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid105]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc105_phy_pc_w))
                begin
                    if(good[long_cpuid105/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid105 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid105/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid105])
        end // if (done[105])

        if (done[106]) begin
            timeout[long_cpuid106] = 0;
            //check_bad_trap(spc106_phy_pc_w, 106, long_cpuid106);
            if(active_thread[long_cpuid106])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc106_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid106/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 106 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid106]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc106_phy_pc_w))
                begin
                    if(good[long_cpuid106/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid106 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid106/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid106])
        end // if (done[106])

        if (done[107]) begin
            timeout[long_cpuid107] = 0;
            //check_bad_trap(spc107_phy_pc_w, 107, long_cpuid107);
            if(active_thread[long_cpuid107])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc107_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid107/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 107 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid107]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc107_phy_pc_w))
                begin
                    if(good[long_cpuid107/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid107 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid107/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid107])
        end // if (done[107])

        if (done[108]) begin
            timeout[long_cpuid108] = 0;
            //check_bad_trap(spc108_phy_pc_w, 108, long_cpuid108);
            if(active_thread[long_cpuid108])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc108_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid108/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 108 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid108]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc108_phy_pc_w))
                begin
                    if(good[long_cpuid108/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid108 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid108/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid108])
        end // if (done[108])

        if (done[109]) begin
            timeout[long_cpuid109] = 0;
            //check_bad_trap(spc109_phy_pc_w, 109, long_cpuid109);
            if(active_thread[long_cpuid109])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc109_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid109/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 109 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid109]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc109_phy_pc_w))
                begin
                    if(good[long_cpuid109/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid109 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid109/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid109])
        end // if (done[109])

        if (done[110]) begin
            timeout[long_cpuid110] = 0;
            //check_bad_trap(spc110_phy_pc_w, 110, long_cpuid110);
            if(active_thread[long_cpuid110])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc110_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid110/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 110 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid110]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc110_phy_pc_w))
                begin
                    if(good[long_cpuid110/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid110 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid110/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid110])
        end // if (done[110])

        if (done[111]) begin
            timeout[long_cpuid111] = 0;
            //check_bad_trap(spc111_phy_pc_w, 111, long_cpuid111);
            if(active_thread[long_cpuid111])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc111_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid111/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 111 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid111]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc111_phy_pc_w))
                begin
                    if(good[long_cpuid111/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid111 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid111/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid111])
        end // if (done[111])

        if (done[112]) begin
            timeout[long_cpuid112] = 0;
            //check_bad_trap(spc112_phy_pc_w, 112, long_cpuid112);
            if(active_thread[long_cpuid112])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc112_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid112/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 112 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid112]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc112_phy_pc_w))
                begin
                    if(good[long_cpuid112/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid112 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid112/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid112])
        end // if (done[112])

        if (done[113]) begin
            timeout[long_cpuid113] = 0;
            //check_bad_trap(spc113_phy_pc_w, 113, long_cpuid113);
            if(active_thread[long_cpuid113])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc113_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid113/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 113 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid113]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc113_phy_pc_w))
                begin
                    if(good[long_cpuid113/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid113 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid113/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid113])
        end // if (done[113])

        if (done[114]) begin
            timeout[long_cpuid114] = 0;
            //check_bad_trap(spc114_phy_pc_w, 114, long_cpuid114);
            if(active_thread[long_cpuid114])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc114_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid114/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 114 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid114]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc114_phy_pc_w))
                begin
                    if(good[long_cpuid114/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid114 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid114/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid114])
        end // if (done[114])

        if (done[115]) begin
            timeout[long_cpuid115] = 0;
            //check_bad_trap(spc115_phy_pc_w, 115, long_cpuid115);
            if(active_thread[long_cpuid115])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc115_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid115/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 115 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid115]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc115_phy_pc_w))
                begin
                    if(good[long_cpuid115/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid115 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid115/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid115])
        end // if (done[115])

        if (done[116]) begin
            timeout[long_cpuid116] = 0;
            //check_bad_trap(spc116_phy_pc_w, 116, long_cpuid116);
            if(active_thread[long_cpuid116])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc116_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid116/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 116 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid116]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc116_phy_pc_w))
                begin
                    if(good[long_cpuid116/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid116 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid116/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid116])
        end // if (done[116])

        if (done[117]) begin
            timeout[long_cpuid117] = 0;
            //check_bad_trap(spc117_phy_pc_w, 117, long_cpuid117);
            if(active_thread[long_cpuid117])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc117_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid117/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 117 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid117]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc117_phy_pc_w))
                begin
                    if(good[long_cpuid117/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid117 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid117/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid117])
        end // if (done[117])

        if (done[118]) begin
            timeout[long_cpuid118] = 0;
            //check_bad_trap(spc118_phy_pc_w, 118, long_cpuid118);
            if(active_thread[long_cpuid118])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc118_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid118/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 118 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid118]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc118_phy_pc_w))
                begin
                    if(good[long_cpuid118/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid118 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid118/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid118])
        end // if (done[118])

        if (done[119]) begin
            timeout[long_cpuid119] = 0;
            //check_bad_trap(spc119_phy_pc_w, 119, long_cpuid119);
            if(active_thread[long_cpuid119])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc119_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid119/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 119 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid119]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc119_phy_pc_w))
                begin
                    if(good[long_cpuid119/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid119 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid119/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid119])
        end // if (done[119])

        if (done[120]) begin
            timeout[long_cpuid120] = 0;
            //check_bad_trap(spc120_phy_pc_w, 120, long_cpuid120);
            if(active_thread[long_cpuid120])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc120_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid120/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 120 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid120]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc120_phy_pc_w))
                begin
                    if(good[long_cpuid120/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid120 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid120/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid120])
        end // if (done[120])

        if (done[121]) begin
            timeout[long_cpuid121] = 0;
            //check_bad_trap(spc121_phy_pc_w, 121, long_cpuid121);
            if(active_thread[long_cpuid121])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc121_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid121/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 121 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid121]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc121_phy_pc_w))
                begin
                    if(good[long_cpuid121/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid121 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid121/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid121])
        end // if (done[121])

        if (done[122]) begin
            timeout[long_cpuid122] = 0;
            //check_bad_trap(spc122_phy_pc_w, 122, long_cpuid122);
            if(active_thread[long_cpuid122])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc122_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid122/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 122 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid122]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc122_phy_pc_w))
                begin
                    if(good[long_cpuid122/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid122 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid122/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid122])
        end // if (done[122])

        if (done[123]) begin
            timeout[long_cpuid123] = 0;
            //check_bad_trap(spc123_phy_pc_w, 123, long_cpuid123);
            if(active_thread[long_cpuid123])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc123_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid123/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 123 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid123]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc123_phy_pc_w))
                begin
                    if(good[long_cpuid123/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid123 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid123/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid123])
        end // if (done[123])

        if (done[124]) begin
            timeout[long_cpuid124] = 0;
            //check_bad_trap(spc124_phy_pc_w, 124, long_cpuid124);
            if(active_thread[long_cpuid124])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc124_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid124/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 124 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid124]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc124_phy_pc_w))
                begin
                    if(good[long_cpuid124/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid124 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid124/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid124])
        end // if (done[124])

        if (done[125]) begin
            timeout[long_cpuid125] = 0;
            //check_bad_trap(spc125_phy_pc_w, 125, long_cpuid125);
            if(active_thread[long_cpuid125])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc125_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid125/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 125 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid125]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc125_phy_pc_w))
                begin
                    if(good[long_cpuid125/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid125 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid125/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid125])
        end // if (done[125])

        if (done[126]) begin
            timeout[long_cpuid126] = 0;
            //check_bad_trap(spc126_phy_pc_w, 126, long_cpuid126);
            if(active_thread[long_cpuid126])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc126_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid126/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 126 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid126]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc126_phy_pc_w))
                begin
                    if(good[long_cpuid126/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid126 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid126/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid126])
        end // if (done[126])

        if (done[127]) begin
            timeout[long_cpuid127] = 0;
            //check_bad_trap(spc127_phy_pc_w, 127, long_cpuid127);
            if(active_thread[long_cpuid127])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc127_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid127/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 127 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid127]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc127_phy_pc_w))
                begin
                    if(good[long_cpuid127/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid127 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid127/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid127])
        end // if (done[127])

        if (done[128]) begin
            timeout[long_cpuid128] = 0;
            //check_bad_trap(spc128_phy_pc_w, 128, long_cpuid128);
            if(active_thread[long_cpuid128])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc128_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid128/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 128 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid128]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc128_phy_pc_w))
                begin
                    if(good[long_cpuid128/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid128 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid128/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid128])
        end // if (done[128])

        if (done[129]) begin
            timeout[long_cpuid129] = 0;
            //check_bad_trap(spc129_phy_pc_w, 129, long_cpuid129);
            if(active_thread[long_cpuid129])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc129_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid129/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 129 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid129]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc129_phy_pc_w))
                begin
                    if(good[long_cpuid129/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid129 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid129/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid129])
        end // if (done[129])

        if (done[130]) begin
            timeout[long_cpuid130] = 0;
            //check_bad_trap(spc130_phy_pc_w, 130, long_cpuid130);
            if(active_thread[long_cpuid130])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc130_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid130/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 130 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid130]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc130_phy_pc_w))
                begin
                    if(good[long_cpuid130/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid130 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid130/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid130])
        end // if (done[130])

        if (done[131]) begin
            timeout[long_cpuid131] = 0;
            //check_bad_trap(spc131_phy_pc_w, 131, long_cpuid131);
            if(active_thread[long_cpuid131])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc131_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid131/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 131 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid131]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc131_phy_pc_w))
                begin
                    if(good[long_cpuid131/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid131 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid131/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid131])
        end // if (done[131])

        if (done[132]) begin
            timeout[long_cpuid132] = 0;
            //check_bad_trap(spc132_phy_pc_w, 132, long_cpuid132);
            if(active_thread[long_cpuid132])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc132_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid132/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 132 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid132]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc132_phy_pc_w))
                begin
                    if(good[long_cpuid132/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid132 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid132/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid132])
        end // if (done[132])

        if (done[133]) begin
            timeout[long_cpuid133] = 0;
            //check_bad_trap(spc133_phy_pc_w, 133, long_cpuid133);
            if(active_thread[long_cpuid133])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc133_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid133/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 133 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid133]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc133_phy_pc_w))
                begin
                    if(good[long_cpuid133/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid133 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid133/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid133])
        end // if (done[133])

        if (done[134]) begin
            timeout[long_cpuid134] = 0;
            //check_bad_trap(spc134_phy_pc_w, 134, long_cpuid134);
            if(active_thread[long_cpuid134])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc134_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid134/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 134 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid134]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc134_phy_pc_w))
                begin
                    if(good[long_cpuid134/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid134 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid134/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid134])
        end // if (done[134])

        if (done[135]) begin
            timeout[long_cpuid135] = 0;
            //check_bad_trap(spc135_phy_pc_w, 135, long_cpuid135);
            if(active_thread[long_cpuid135])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc135_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid135/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 135 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid135]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc135_phy_pc_w))
                begin
                    if(good[long_cpuid135/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid135 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid135/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid135])
        end // if (done[135])

        if (done[136]) begin
            timeout[long_cpuid136] = 0;
            //check_bad_trap(spc136_phy_pc_w, 136, long_cpuid136);
            if(active_thread[long_cpuid136])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc136_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid136/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 136 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid136]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc136_phy_pc_w))
                begin
                    if(good[long_cpuid136/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid136 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid136/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid136])
        end // if (done[136])

        if (done[137]) begin
            timeout[long_cpuid137] = 0;
            //check_bad_trap(spc137_phy_pc_w, 137, long_cpuid137);
            if(active_thread[long_cpuid137])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc137_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid137/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 137 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid137]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc137_phy_pc_w))
                begin
                    if(good[long_cpuid137/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid137 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid137/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid137])
        end // if (done[137])

        if (done[138]) begin
            timeout[long_cpuid138] = 0;
            //check_bad_trap(spc138_phy_pc_w, 138, long_cpuid138);
            if(active_thread[long_cpuid138])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc138_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid138/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 138 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid138]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc138_phy_pc_w))
                begin
                    if(good[long_cpuid138/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid138 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid138/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid138])
        end // if (done[138])

        if (done[139]) begin
            timeout[long_cpuid139] = 0;
            //check_bad_trap(spc139_phy_pc_w, 139, long_cpuid139);
            if(active_thread[long_cpuid139])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc139_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid139/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 139 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid139]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc139_phy_pc_w))
                begin
                    if(good[long_cpuid139/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid139 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid139/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid139])
        end // if (done[139])

        if (done[140]) begin
            timeout[long_cpuid140] = 0;
            //check_bad_trap(spc140_phy_pc_w, 140, long_cpuid140);
            if(active_thread[long_cpuid140])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc140_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid140/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 140 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid140]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc140_phy_pc_w))
                begin
                    if(good[long_cpuid140/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid140 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid140/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid140])
        end // if (done[140])

        if (done[141]) begin
            timeout[long_cpuid141] = 0;
            //check_bad_trap(spc141_phy_pc_w, 141, long_cpuid141);
            if(active_thread[long_cpuid141])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc141_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid141/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 141 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid141]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc141_phy_pc_w))
                begin
                    if(good[long_cpuid141/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid141 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid141/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid141])
        end // if (done[141])

        if (done[142]) begin
            timeout[long_cpuid142] = 0;
            //check_bad_trap(spc142_phy_pc_w, 142, long_cpuid142);
            if(active_thread[long_cpuid142])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc142_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid142/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 142 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid142]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc142_phy_pc_w))
                begin
                    if(good[long_cpuid142/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid142 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid142/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid142])
        end // if (done[142])

        if (done[143]) begin
            timeout[long_cpuid143] = 0;
            //check_bad_trap(spc143_phy_pc_w, 143, long_cpuid143);
            if(active_thread[long_cpuid143])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc143_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid143/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 143 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid143]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc143_phy_pc_w))
                begin
                    if(good[long_cpuid143/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid143 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid143/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid143])
        end // if (done[143])

        if (done[144]) begin
            timeout[long_cpuid144] = 0;
            //check_bad_trap(spc144_phy_pc_w, 144, long_cpuid144);
            if(active_thread[long_cpuid144])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc144_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid144/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 144 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid144]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc144_phy_pc_w))
                begin
                    if(good[long_cpuid144/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid144 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid144/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid144])
        end // if (done[144])

        if (done[145]) begin
            timeout[long_cpuid145] = 0;
            //check_bad_trap(spc145_phy_pc_w, 145, long_cpuid145);
            if(active_thread[long_cpuid145])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc145_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid145/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 145 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid145]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc145_phy_pc_w))
                begin
                    if(good[long_cpuid145/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid145 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid145/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid145])
        end // if (done[145])

        if (done[146]) begin
            timeout[long_cpuid146] = 0;
            //check_bad_trap(spc146_phy_pc_w, 146, long_cpuid146);
            if(active_thread[long_cpuid146])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc146_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid146/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 146 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid146]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc146_phy_pc_w))
                begin
                    if(good[long_cpuid146/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid146 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid146/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid146])
        end // if (done[146])

        if (done[147]) begin
            timeout[long_cpuid147] = 0;
            //check_bad_trap(spc147_phy_pc_w, 147, long_cpuid147);
            if(active_thread[long_cpuid147])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc147_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid147/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 147 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid147]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc147_phy_pc_w))
                begin
                    if(good[long_cpuid147/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid147 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid147/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid147])
        end // if (done[147])

        if (done[148]) begin
            timeout[long_cpuid148] = 0;
            //check_bad_trap(spc148_phy_pc_w, 148, long_cpuid148);
            if(active_thread[long_cpuid148])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc148_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid148/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 148 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid148]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc148_phy_pc_w))
                begin
                    if(good[long_cpuid148/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid148 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid148/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid148])
        end // if (done[148])

        if (done[149]) begin
            timeout[long_cpuid149] = 0;
            //check_bad_trap(spc149_phy_pc_w, 149, long_cpuid149);
            if(active_thread[long_cpuid149])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc149_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid149/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 149 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid149]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc149_phy_pc_w))
                begin
                    if(good[long_cpuid149/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid149 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid149/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid149])
        end // if (done[149])

        if (done[150]) begin
            timeout[long_cpuid150] = 0;
            //check_bad_trap(spc150_phy_pc_w, 150, long_cpuid150);
            if(active_thread[long_cpuid150])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc150_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid150/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 150 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid150]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc150_phy_pc_w))
                begin
                    if(good[long_cpuid150/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid150 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid150/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid150])
        end // if (done[150])

        if (done[151]) begin
            timeout[long_cpuid151] = 0;
            //check_bad_trap(spc151_phy_pc_w, 151, long_cpuid151);
            if(active_thread[long_cpuid151])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc151_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid151/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 151 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid151]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc151_phy_pc_w))
                begin
                    if(good[long_cpuid151/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid151 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid151/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid151])
        end // if (done[151])

        if (done[152]) begin
            timeout[long_cpuid152] = 0;
            //check_bad_trap(spc152_phy_pc_w, 152, long_cpuid152);
            if(active_thread[long_cpuid152])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc152_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid152/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 152 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid152]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc152_phy_pc_w))
                begin
                    if(good[long_cpuid152/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid152 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid152/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid152])
        end // if (done[152])

        if (done[153]) begin
            timeout[long_cpuid153] = 0;
            //check_bad_trap(spc153_phy_pc_w, 153, long_cpuid153);
            if(active_thread[long_cpuid153])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc153_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid153/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 153 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid153]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc153_phy_pc_w))
                begin
                    if(good[long_cpuid153/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid153 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid153/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid153])
        end // if (done[153])

        if (done[154]) begin
            timeout[long_cpuid154] = 0;
            //check_bad_trap(spc154_phy_pc_w, 154, long_cpuid154);
            if(active_thread[long_cpuid154])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc154_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid154/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 154 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid154]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc154_phy_pc_w))
                begin
                    if(good[long_cpuid154/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid154 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid154/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid154])
        end // if (done[154])

        if (done[155]) begin
            timeout[long_cpuid155] = 0;
            //check_bad_trap(spc155_phy_pc_w, 155, long_cpuid155);
            if(active_thread[long_cpuid155])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc155_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid155/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 155 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid155]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc155_phy_pc_w))
                begin
                    if(good[long_cpuid155/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid155 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid155/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid155])
        end // if (done[155])

        if (done[156]) begin
            timeout[long_cpuid156] = 0;
            //check_bad_trap(spc156_phy_pc_w, 156, long_cpuid156);
            if(active_thread[long_cpuid156])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc156_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid156/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 156 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid156]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc156_phy_pc_w))
                begin
                    if(good[long_cpuid156/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid156 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid156/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid156])
        end // if (done[156])

        if (done[157]) begin
            timeout[long_cpuid157] = 0;
            //check_bad_trap(spc157_phy_pc_w, 157, long_cpuid157);
            if(active_thread[long_cpuid157])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc157_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid157/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 157 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid157]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc157_phy_pc_w))
                begin
                    if(good[long_cpuid157/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid157 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid157/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid157])
        end // if (done[157])

        if (done[158]) begin
            timeout[long_cpuid158] = 0;
            //check_bad_trap(spc158_phy_pc_w, 158, long_cpuid158);
            if(active_thread[long_cpuid158])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc158_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid158/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 158 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid158]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc158_phy_pc_w))
                begin
                    if(good[long_cpuid158/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid158 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid158/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid158])
        end // if (done[158])

        if (done[159]) begin
            timeout[long_cpuid159] = 0;
            //check_bad_trap(spc159_phy_pc_w, 159, long_cpuid159);
            if(active_thread[long_cpuid159])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc159_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid159/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 159 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid159]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc159_phy_pc_w))
                begin
                    if(good[long_cpuid159/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid159 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid159/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid159])
        end // if (done[159])

        if (done[160]) begin
            timeout[long_cpuid160] = 0;
            //check_bad_trap(spc160_phy_pc_w, 160, long_cpuid160);
            if(active_thread[long_cpuid160])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc160_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid160/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 160 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid160]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc160_phy_pc_w))
                begin
                    if(good[long_cpuid160/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid160 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid160/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid160])
        end // if (done[160])

        if (done[161]) begin
            timeout[long_cpuid161] = 0;
            //check_bad_trap(spc161_phy_pc_w, 161, long_cpuid161);
            if(active_thread[long_cpuid161])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc161_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid161/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 161 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid161]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc161_phy_pc_w))
                begin
                    if(good[long_cpuid161/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid161 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid161/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid161])
        end // if (done[161])

        if (done[162]) begin
            timeout[long_cpuid162] = 0;
            //check_bad_trap(spc162_phy_pc_w, 162, long_cpuid162);
            if(active_thread[long_cpuid162])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc162_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid162/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 162 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid162]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc162_phy_pc_w))
                begin
                    if(good[long_cpuid162/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid162 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid162/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid162])
        end // if (done[162])

        if (done[163]) begin
            timeout[long_cpuid163] = 0;
            //check_bad_trap(spc163_phy_pc_w, 163, long_cpuid163);
            if(active_thread[long_cpuid163])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc163_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid163/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 163 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid163]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc163_phy_pc_w))
                begin
                    if(good[long_cpuid163/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid163 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid163/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid163])
        end // if (done[163])

        if (done[164]) begin
            timeout[long_cpuid164] = 0;
            //check_bad_trap(spc164_phy_pc_w, 164, long_cpuid164);
            if(active_thread[long_cpuid164])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc164_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid164/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 164 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid164]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc164_phy_pc_w))
                begin
                    if(good[long_cpuid164/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid164 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid164/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid164])
        end // if (done[164])

        if (done[165]) begin
            timeout[long_cpuid165] = 0;
            //check_bad_trap(spc165_phy_pc_w, 165, long_cpuid165);
            if(active_thread[long_cpuid165])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc165_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid165/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 165 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid165]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc165_phy_pc_w))
                begin
                    if(good[long_cpuid165/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid165 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid165/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid165])
        end // if (done[165])

        if (done[166]) begin
            timeout[long_cpuid166] = 0;
            //check_bad_trap(spc166_phy_pc_w, 166, long_cpuid166);
            if(active_thread[long_cpuid166])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc166_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid166/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 166 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid166]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc166_phy_pc_w))
                begin
                    if(good[long_cpuid166/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid166 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid166/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid166])
        end // if (done[166])

        if (done[167]) begin
            timeout[long_cpuid167] = 0;
            //check_bad_trap(spc167_phy_pc_w, 167, long_cpuid167);
            if(active_thread[long_cpuid167])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc167_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid167/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 167 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid167]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc167_phy_pc_w))
                begin
                    if(good[long_cpuid167/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid167 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid167/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid167])
        end // if (done[167])

        if (done[168]) begin
            timeout[long_cpuid168] = 0;
            //check_bad_trap(spc168_phy_pc_w, 168, long_cpuid168);
            if(active_thread[long_cpuid168])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc168_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid168/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 168 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid168]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc168_phy_pc_w))
                begin
                    if(good[long_cpuid168/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid168 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid168/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid168])
        end // if (done[168])

        if (done[169]) begin
            timeout[long_cpuid169] = 0;
            //check_bad_trap(spc169_phy_pc_w, 169, long_cpuid169);
            if(active_thread[long_cpuid169])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc169_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid169/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 169 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid169]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc169_phy_pc_w))
                begin
                    if(good[long_cpuid169/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid169 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid169/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid169])
        end // if (done[169])

        if (done[170]) begin
            timeout[long_cpuid170] = 0;
            //check_bad_trap(spc170_phy_pc_w, 170, long_cpuid170);
            if(active_thread[long_cpuid170])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc170_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid170/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 170 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid170]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc170_phy_pc_w))
                begin
                    if(good[long_cpuid170/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid170 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid170/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid170])
        end // if (done[170])

        if (done[171]) begin
            timeout[long_cpuid171] = 0;
            //check_bad_trap(spc171_phy_pc_w, 171, long_cpuid171);
            if(active_thread[long_cpuid171])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc171_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid171/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 171 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid171]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc171_phy_pc_w))
                begin
                    if(good[long_cpuid171/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid171 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid171/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid171])
        end // if (done[171])

        if (done[172]) begin
            timeout[long_cpuid172] = 0;
            //check_bad_trap(spc172_phy_pc_w, 172, long_cpuid172);
            if(active_thread[long_cpuid172])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc172_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid172/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 172 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid172]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc172_phy_pc_w))
                begin
                    if(good[long_cpuid172/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid172 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid172/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid172])
        end // if (done[172])

        if (done[173]) begin
            timeout[long_cpuid173] = 0;
            //check_bad_trap(spc173_phy_pc_w, 173, long_cpuid173);
            if(active_thread[long_cpuid173])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc173_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid173/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 173 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid173]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc173_phy_pc_w))
                begin
                    if(good[long_cpuid173/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid173 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid173/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid173])
        end // if (done[173])

        if (done[174]) begin
            timeout[long_cpuid174] = 0;
            //check_bad_trap(spc174_phy_pc_w, 174, long_cpuid174);
            if(active_thread[long_cpuid174])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc174_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid174/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 174 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid174]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc174_phy_pc_w))
                begin
                    if(good[long_cpuid174/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid174 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid174/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid174])
        end // if (done[174])

        if (done[175]) begin
            timeout[long_cpuid175] = 0;
            //check_bad_trap(spc175_phy_pc_w, 175, long_cpuid175);
            if(active_thread[long_cpuid175])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc175_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid175/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 175 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid175]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc175_phy_pc_w))
                begin
                    if(good[long_cpuid175/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid175 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid175/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid175])
        end // if (done[175])

        if (done[176]) begin
            timeout[long_cpuid176] = 0;
            //check_bad_trap(spc176_phy_pc_w, 176, long_cpuid176);
            if(active_thread[long_cpuid176])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc176_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid176/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 176 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid176]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc176_phy_pc_w))
                begin
                    if(good[long_cpuid176/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid176 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid176/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid176])
        end // if (done[176])

        if (done[177]) begin
            timeout[long_cpuid177] = 0;
            //check_bad_trap(spc177_phy_pc_w, 177, long_cpuid177);
            if(active_thread[long_cpuid177])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc177_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid177/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 177 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid177]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc177_phy_pc_w))
                begin
                    if(good[long_cpuid177/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid177 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid177/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid177])
        end // if (done[177])

        if (done[178]) begin
            timeout[long_cpuid178] = 0;
            //check_bad_trap(spc178_phy_pc_w, 178, long_cpuid178);
            if(active_thread[long_cpuid178])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc178_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid178/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 178 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid178]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc178_phy_pc_w))
                begin
                    if(good[long_cpuid178/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid178 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid178/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid178])
        end // if (done[178])

        if (done[179]) begin
            timeout[long_cpuid179] = 0;
            //check_bad_trap(spc179_phy_pc_w, 179, long_cpuid179);
            if(active_thread[long_cpuid179])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc179_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid179/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 179 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid179]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc179_phy_pc_w))
                begin
                    if(good[long_cpuid179/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid179 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid179/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid179])
        end // if (done[179])

        if (done[180]) begin
            timeout[long_cpuid180] = 0;
            //check_bad_trap(spc180_phy_pc_w, 180, long_cpuid180);
            if(active_thread[long_cpuid180])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc180_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid180/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 180 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid180]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc180_phy_pc_w))
                begin
                    if(good[long_cpuid180/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid180 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid180/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid180])
        end // if (done[180])

        if (done[181]) begin
            timeout[long_cpuid181] = 0;
            //check_bad_trap(spc181_phy_pc_w, 181, long_cpuid181);
            if(active_thread[long_cpuid181])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc181_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid181/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 181 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid181]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc181_phy_pc_w))
                begin
                    if(good[long_cpuid181/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid181 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid181/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid181])
        end // if (done[181])

        if (done[182]) begin
            timeout[long_cpuid182] = 0;
            //check_bad_trap(spc182_phy_pc_w, 182, long_cpuid182);
            if(active_thread[long_cpuid182])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc182_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid182/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 182 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid182]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc182_phy_pc_w))
                begin
                    if(good[long_cpuid182/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid182 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid182/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid182])
        end // if (done[182])

        if (done[183]) begin
            timeout[long_cpuid183] = 0;
            //check_bad_trap(spc183_phy_pc_w, 183, long_cpuid183);
            if(active_thread[long_cpuid183])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc183_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid183/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 183 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid183]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc183_phy_pc_w))
                begin
                    if(good[long_cpuid183/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid183 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid183/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid183])
        end // if (done[183])

        if (done[184]) begin
            timeout[long_cpuid184] = 0;
            //check_bad_trap(spc184_phy_pc_w, 184, long_cpuid184);
            if(active_thread[long_cpuid184])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc184_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid184/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 184 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid184]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc184_phy_pc_w))
                begin
                    if(good[long_cpuid184/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid184 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid184/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid184])
        end // if (done[184])

        if (done[185]) begin
            timeout[long_cpuid185] = 0;
            //check_bad_trap(spc185_phy_pc_w, 185, long_cpuid185);
            if(active_thread[long_cpuid185])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc185_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid185/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 185 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid185]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc185_phy_pc_w))
                begin
                    if(good[long_cpuid185/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid185 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid185/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid185])
        end // if (done[185])

        if (done[186]) begin
            timeout[long_cpuid186] = 0;
            //check_bad_trap(spc186_phy_pc_w, 186, long_cpuid186);
            if(active_thread[long_cpuid186])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc186_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid186/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 186 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid186]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc186_phy_pc_w))
                begin
                    if(good[long_cpuid186/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid186 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid186/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid186])
        end // if (done[186])

        if (done[187]) begin
            timeout[long_cpuid187] = 0;
            //check_bad_trap(spc187_phy_pc_w, 187, long_cpuid187);
            if(active_thread[long_cpuid187])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc187_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid187/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 187 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid187]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc187_phy_pc_w))
                begin
                    if(good[long_cpuid187/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid187 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid187/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid187])
        end // if (done[187])

        if (done[188]) begin
            timeout[long_cpuid188] = 0;
            //check_bad_trap(spc188_phy_pc_w, 188, long_cpuid188);
            if(active_thread[long_cpuid188])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc188_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid188/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 188 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid188]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc188_phy_pc_w))
                begin
                    if(good[long_cpuid188/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid188 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid188/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid188])
        end // if (done[188])

        if (done[189]) begin
            timeout[long_cpuid189] = 0;
            //check_bad_trap(spc189_phy_pc_w, 189, long_cpuid189);
            if(active_thread[long_cpuid189])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc189_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid189/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 189 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid189]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc189_phy_pc_w))
                begin
                    if(good[long_cpuid189/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid189 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid189/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid189])
        end // if (done[189])

        if (done[190]) begin
            timeout[long_cpuid190] = 0;
            //check_bad_trap(spc190_phy_pc_w, 190, long_cpuid190);
            if(active_thread[long_cpuid190])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc190_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid190/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 190 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid190]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc190_phy_pc_w))
                begin
                    if(good[long_cpuid190/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid190 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid190/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid190])
        end // if (done[190])

        if (done[191]) begin
            timeout[long_cpuid191] = 0;
            //check_bad_trap(spc191_phy_pc_w, 191, long_cpuid191);
            if(active_thread[long_cpuid191])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc191_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid191/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 191 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid191]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc191_phy_pc_w))
                begin
                    if(good[long_cpuid191/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid191 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid191/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid191])
        end // if (done[191])

        if (done[192]) begin
            timeout[long_cpuid192] = 0;
            //check_bad_trap(spc192_phy_pc_w, 192, long_cpuid192);
            if(active_thread[long_cpuid192])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc192_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid192/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 192 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid192]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc192_phy_pc_w))
                begin
                    if(good[long_cpuid192/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid192 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid192/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid192])
        end // if (done[192])

        if (done[193]) begin
            timeout[long_cpuid193] = 0;
            //check_bad_trap(spc193_phy_pc_w, 193, long_cpuid193);
            if(active_thread[long_cpuid193])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc193_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid193/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 193 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid193]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc193_phy_pc_w))
                begin
                    if(good[long_cpuid193/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid193 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid193/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid193])
        end // if (done[193])

        if (done[194]) begin
            timeout[long_cpuid194] = 0;
            //check_bad_trap(spc194_phy_pc_w, 194, long_cpuid194);
            if(active_thread[long_cpuid194])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc194_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid194/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 194 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid194]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc194_phy_pc_w))
                begin
                    if(good[long_cpuid194/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid194 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid194/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid194])
        end // if (done[194])

        if (done[195]) begin
            timeout[long_cpuid195] = 0;
            //check_bad_trap(spc195_phy_pc_w, 195, long_cpuid195);
            if(active_thread[long_cpuid195])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc195_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid195/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 195 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid195]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc195_phy_pc_w))
                begin
                    if(good[long_cpuid195/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid195 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid195/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid195])
        end // if (done[195])

        if (done[196]) begin
            timeout[long_cpuid196] = 0;
            //check_bad_trap(spc196_phy_pc_w, 196, long_cpuid196);
            if(active_thread[long_cpuid196])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc196_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid196/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 196 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid196]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc196_phy_pc_w))
                begin
                    if(good[long_cpuid196/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid196 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid196/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid196])
        end // if (done[196])

        if (done[197]) begin
            timeout[long_cpuid197] = 0;
            //check_bad_trap(spc197_phy_pc_w, 197, long_cpuid197);
            if(active_thread[long_cpuid197])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc197_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid197/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 197 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid197]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc197_phy_pc_w))
                begin
                    if(good[long_cpuid197/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid197 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid197/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid197])
        end // if (done[197])

        if (done[198]) begin
            timeout[long_cpuid198] = 0;
            //check_bad_trap(spc198_phy_pc_w, 198, long_cpuid198);
            if(active_thread[long_cpuid198])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc198_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid198/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 198 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid198]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc198_phy_pc_w))
                begin
                    if(good[long_cpuid198/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid198 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid198/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid198])
        end // if (done[198])

        if (done[199]) begin
            timeout[long_cpuid199] = 0;
            //check_bad_trap(spc199_phy_pc_w, 199, long_cpuid199);
            if(active_thread[long_cpuid199])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc199_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid199/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 199 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid199]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc199_phy_pc_w))
                begin
                    if(good[long_cpuid199/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid199 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid199/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid199])
        end // if (done[199])

        if (done[200]) begin
            timeout[long_cpuid200] = 0;
            //check_bad_trap(spc200_phy_pc_w, 200, long_cpuid200);
            if(active_thread[long_cpuid200])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc200_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid200/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 200 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid200]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc200_phy_pc_w))
                begin
                    if(good[long_cpuid200/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid200 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid200/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid200])
        end // if (done[200])

        if (done[201]) begin
            timeout[long_cpuid201] = 0;
            //check_bad_trap(spc201_phy_pc_w, 201, long_cpuid201);
            if(active_thread[long_cpuid201])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc201_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid201/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 201 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid201]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc201_phy_pc_w))
                begin
                    if(good[long_cpuid201/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid201 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid201/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid201])
        end // if (done[201])

        if (done[202]) begin
            timeout[long_cpuid202] = 0;
            //check_bad_trap(spc202_phy_pc_w, 202, long_cpuid202);
            if(active_thread[long_cpuid202])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc202_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid202/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 202 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid202]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc202_phy_pc_w))
                begin
                    if(good[long_cpuid202/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid202 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid202/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid202])
        end // if (done[202])

        if (done[203]) begin
            timeout[long_cpuid203] = 0;
            //check_bad_trap(spc203_phy_pc_w, 203, long_cpuid203);
            if(active_thread[long_cpuid203])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc203_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid203/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 203 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid203]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc203_phy_pc_w))
                begin
                    if(good[long_cpuid203/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid203 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid203/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid203])
        end // if (done[203])

        if (done[204]) begin
            timeout[long_cpuid204] = 0;
            //check_bad_trap(spc204_phy_pc_w, 204, long_cpuid204);
            if(active_thread[long_cpuid204])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc204_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid204/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 204 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid204]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc204_phy_pc_w))
                begin
                    if(good[long_cpuid204/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid204 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid204/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid204])
        end // if (done[204])

        if (done[205]) begin
            timeout[long_cpuid205] = 0;
            //check_bad_trap(spc205_phy_pc_w, 205, long_cpuid205);
            if(active_thread[long_cpuid205])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc205_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid205/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 205 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid205]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc205_phy_pc_w))
                begin
                    if(good[long_cpuid205/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid205 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid205/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid205])
        end // if (done[205])

        if (done[206]) begin
            timeout[long_cpuid206] = 0;
            //check_bad_trap(spc206_phy_pc_w, 206, long_cpuid206);
            if(active_thread[long_cpuid206])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc206_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid206/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 206 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid206]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc206_phy_pc_w))
                begin
                    if(good[long_cpuid206/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid206 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid206/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid206])
        end // if (done[206])

        if (done[207]) begin
            timeout[long_cpuid207] = 0;
            //check_bad_trap(spc207_phy_pc_w, 207, long_cpuid207);
            if(active_thread[long_cpuid207])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc207_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid207/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 207 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid207]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc207_phy_pc_w))
                begin
                    if(good[long_cpuid207/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid207 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid207/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid207])
        end // if (done[207])

        if (done[208]) begin
            timeout[long_cpuid208] = 0;
            //check_bad_trap(spc208_phy_pc_w, 208, long_cpuid208);
            if(active_thread[long_cpuid208])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc208_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid208/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 208 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid208]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc208_phy_pc_w))
                begin
                    if(good[long_cpuid208/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid208 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid208/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid208])
        end // if (done[208])

        if (done[209]) begin
            timeout[long_cpuid209] = 0;
            //check_bad_trap(spc209_phy_pc_w, 209, long_cpuid209);
            if(active_thread[long_cpuid209])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc209_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid209/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 209 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid209]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc209_phy_pc_w))
                begin
                    if(good[long_cpuid209/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid209 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid209/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid209])
        end // if (done[209])

        if (done[210]) begin
            timeout[long_cpuid210] = 0;
            //check_bad_trap(spc210_phy_pc_w, 210, long_cpuid210);
            if(active_thread[long_cpuid210])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc210_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid210/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 210 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid210]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc210_phy_pc_w))
                begin
                    if(good[long_cpuid210/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid210 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid210/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid210])
        end // if (done[210])

        if (done[211]) begin
            timeout[long_cpuid211] = 0;
            //check_bad_trap(spc211_phy_pc_w, 211, long_cpuid211);
            if(active_thread[long_cpuid211])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc211_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid211/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 211 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid211]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc211_phy_pc_w))
                begin
                    if(good[long_cpuid211/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid211 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid211/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid211])
        end // if (done[211])

        if (done[212]) begin
            timeout[long_cpuid212] = 0;
            //check_bad_trap(spc212_phy_pc_w, 212, long_cpuid212);
            if(active_thread[long_cpuid212])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc212_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid212/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 212 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid212]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc212_phy_pc_w))
                begin
                    if(good[long_cpuid212/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid212 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid212/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid212])
        end // if (done[212])

        if (done[213]) begin
            timeout[long_cpuid213] = 0;
            //check_bad_trap(spc213_phy_pc_w, 213, long_cpuid213);
            if(active_thread[long_cpuid213])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc213_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid213/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 213 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid213]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc213_phy_pc_w))
                begin
                    if(good[long_cpuid213/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid213 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid213/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid213])
        end // if (done[213])

        if (done[214]) begin
            timeout[long_cpuid214] = 0;
            //check_bad_trap(spc214_phy_pc_w, 214, long_cpuid214);
            if(active_thread[long_cpuid214])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc214_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid214/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 214 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid214]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc214_phy_pc_w))
                begin
                    if(good[long_cpuid214/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid214 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid214/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid214])
        end // if (done[214])

        if (done[215]) begin
            timeout[long_cpuid215] = 0;
            //check_bad_trap(spc215_phy_pc_w, 215, long_cpuid215);
            if(active_thread[long_cpuid215])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc215_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid215/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 215 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid215]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc215_phy_pc_w))
                begin
                    if(good[long_cpuid215/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid215 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid215/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid215])
        end // if (done[215])

        if (done[216]) begin
            timeout[long_cpuid216] = 0;
            //check_bad_trap(spc216_phy_pc_w, 216, long_cpuid216);
            if(active_thread[long_cpuid216])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc216_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid216/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 216 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid216]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc216_phy_pc_w))
                begin
                    if(good[long_cpuid216/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid216 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid216/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid216])
        end // if (done[216])

        if (done[217]) begin
            timeout[long_cpuid217] = 0;
            //check_bad_trap(spc217_phy_pc_w, 217, long_cpuid217);
            if(active_thread[long_cpuid217])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc217_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid217/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 217 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid217]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc217_phy_pc_w))
                begin
                    if(good[long_cpuid217/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid217 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid217/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid217])
        end // if (done[217])

        if (done[218]) begin
            timeout[long_cpuid218] = 0;
            //check_bad_trap(spc218_phy_pc_w, 218, long_cpuid218);
            if(active_thread[long_cpuid218])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc218_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid218/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 218 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid218]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc218_phy_pc_w))
                begin
                    if(good[long_cpuid218/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid218 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid218/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid218])
        end // if (done[218])

        if (done[219]) begin
            timeout[long_cpuid219] = 0;
            //check_bad_trap(spc219_phy_pc_w, 219, long_cpuid219);
            if(active_thread[long_cpuid219])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc219_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid219/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 219 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid219]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc219_phy_pc_w))
                begin
                    if(good[long_cpuid219/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid219 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid219/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid219])
        end // if (done[219])

        if (done[220]) begin
            timeout[long_cpuid220] = 0;
            //check_bad_trap(spc220_phy_pc_w, 220, long_cpuid220);
            if(active_thread[long_cpuid220])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc220_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid220/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 220 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid220]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc220_phy_pc_w))
                begin
                    if(good[long_cpuid220/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid220 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid220/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid220])
        end // if (done[220])

        if (done[221]) begin
            timeout[long_cpuid221] = 0;
            //check_bad_trap(spc221_phy_pc_w, 221, long_cpuid221);
            if(active_thread[long_cpuid221])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc221_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid221/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 221 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid221]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc221_phy_pc_w))
                begin
                    if(good[long_cpuid221/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid221 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid221/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid221])
        end // if (done[221])

        if (done[222]) begin
            timeout[long_cpuid222] = 0;
            //check_bad_trap(spc222_phy_pc_w, 222, long_cpuid222);
            if(active_thread[long_cpuid222])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc222_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid222/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 222 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid222]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc222_phy_pc_w))
                begin
                    if(good[long_cpuid222/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid222 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid222/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid222])
        end // if (done[222])

        if (done[223]) begin
            timeout[long_cpuid223] = 0;
            //check_bad_trap(spc223_phy_pc_w, 223, long_cpuid223);
            if(active_thread[long_cpuid223])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc223_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid223/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 223 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid223]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc223_phy_pc_w))
                begin
                    if(good[long_cpuid223/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid223 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid223/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid223])
        end // if (done[223])

        if (done[224]) begin
            timeout[long_cpuid224] = 0;
            //check_bad_trap(spc224_phy_pc_w, 224, long_cpuid224);
            if(active_thread[long_cpuid224])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc224_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid224/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 224 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid224]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc224_phy_pc_w))
                begin
                    if(good[long_cpuid224/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid224 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid224/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid224])
        end // if (done[224])

        if (done[225]) begin
            timeout[long_cpuid225] = 0;
            //check_bad_trap(spc225_phy_pc_w, 225, long_cpuid225);
            if(active_thread[long_cpuid225])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc225_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid225/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 225 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid225]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc225_phy_pc_w))
                begin
                    if(good[long_cpuid225/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid225 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid225/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid225])
        end // if (done[225])

        if (done[226]) begin
            timeout[long_cpuid226] = 0;
            //check_bad_trap(spc226_phy_pc_w, 226, long_cpuid226);
            if(active_thread[long_cpuid226])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc226_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid226/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 226 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid226]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc226_phy_pc_w))
                begin
                    if(good[long_cpuid226/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid226 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid226/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid226])
        end // if (done[226])

        if (done[227]) begin
            timeout[long_cpuid227] = 0;
            //check_bad_trap(spc227_phy_pc_w, 227, long_cpuid227);
            if(active_thread[long_cpuid227])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc227_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid227/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 227 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid227]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc227_phy_pc_w))
                begin
                    if(good[long_cpuid227/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid227 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid227/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid227])
        end // if (done[227])

        if (done[228]) begin
            timeout[long_cpuid228] = 0;
            //check_bad_trap(spc228_phy_pc_w, 228, long_cpuid228);
            if(active_thread[long_cpuid228])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc228_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid228/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 228 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid228]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc228_phy_pc_w))
                begin
                    if(good[long_cpuid228/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid228 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid228/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid228])
        end // if (done[228])

        if (done[229]) begin
            timeout[long_cpuid229] = 0;
            //check_bad_trap(spc229_phy_pc_w, 229, long_cpuid229);
            if(active_thread[long_cpuid229])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc229_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid229/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 229 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid229]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc229_phy_pc_w))
                begin
                    if(good[long_cpuid229/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid229 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid229/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid229])
        end // if (done[229])

        if (done[230]) begin
            timeout[long_cpuid230] = 0;
            //check_bad_trap(spc230_phy_pc_w, 230, long_cpuid230);
            if(active_thread[long_cpuid230])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc230_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid230/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 230 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid230]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc230_phy_pc_w))
                begin
                    if(good[long_cpuid230/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid230 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid230/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid230])
        end // if (done[230])

        if (done[231]) begin
            timeout[long_cpuid231] = 0;
            //check_bad_trap(spc231_phy_pc_w, 231, long_cpuid231);
            if(active_thread[long_cpuid231])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc231_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid231/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 231 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid231]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc231_phy_pc_w))
                begin
                    if(good[long_cpuid231/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid231 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid231/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid231])
        end // if (done[231])

        if (done[232]) begin
            timeout[long_cpuid232] = 0;
            //check_bad_trap(spc232_phy_pc_w, 232, long_cpuid232);
            if(active_thread[long_cpuid232])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc232_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid232/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 232 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid232]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc232_phy_pc_w))
                begin
                    if(good[long_cpuid232/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid232 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid232/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid232])
        end // if (done[232])

        if (done[233]) begin
            timeout[long_cpuid233] = 0;
            //check_bad_trap(spc233_phy_pc_w, 233, long_cpuid233);
            if(active_thread[long_cpuid233])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc233_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid233/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 233 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid233]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc233_phy_pc_w))
                begin
                    if(good[long_cpuid233/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid233 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid233/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid233])
        end // if (done[233])

        if (done[234]) begin
            timeout[long_cpuid234] = 0;
            //check_bad_trap(spc234_phy_pc_w, 234, long_cpuid234);
            if(active_thread[long_cpuid234])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc234_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid234/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 234 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid234]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc234_phy_pc_w))
                begin
                    if(good[long_cpuid234/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid234 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid234/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid234])
        end // if (done[234])

        if (done[235]) begin
            timeout[long_cpuid235] = 0;
            //check_bad_trap(spc235_phy_pc_w, 235, long_cpuid235);
            if(active_thread[long_cpuid235])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc235_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid235/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 235 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid235]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc235_phy_pc_w))
                begin
                    if(good[long_cpuid235/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid235 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid235/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid235])
        end // if (done[235])

        if (done[236]) begin
            timeout[long_cpuid236] = 0;
            //check_bad_trap(spc236_phy_pc_w, 236, long_cpuid236);
            if(active_thread[long_cpuid236])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc236_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid236/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 236 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid236]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc236_phy_pc_w))
                begin
                    if(good[long_cpuid236/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid236 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid236/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid236])
        end // if (done[236])

        if (done[237]) begin
            timeout[long_cpuid237] = 0;
            //check_bad_trap(spc237_phy_pc_w, 237, long_cpuid237);
            if(active_thread[long_cpuid237])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc237_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid237/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 237 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid237]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc237_phy_pc_w))
                begin
                    if(good[long_cpuid237/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid237 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid237/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid237])
        end // if (done[237])

        if (done[238]) begin
            timeout[long_cpuid238] = 0;
            //check_bad_trap(spc238_phy_pc_w, 238, long_cpuid238);
            if(active_thread[long_cpuid238])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc238_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid238/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 238 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid238]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc238_phy_pc_w))
                begin
                    if(good[long_cpuid238/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid238 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid238/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid238])
        end // if (done[238])

        if (done[239]) begin
            timeout[long_cpuid239] = 0;
            //check_bad_trap(spc239_phy_pc_w, 239, long_cpuid239);
            if(active_thread[long_cpuid239])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc239_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid239/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 239 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid239]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc239_phy_pc_w))
                begin
                    if(good[long_cpuid239/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid239 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid239/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid239])
        end // if (done[239])

        if (done[240]) begin
            timeout[long_cpuid240] = 0;
            //check_bad_trap(spc240_phy_pc_w, 240, long_cpuid240);
            if(active_thread[long_cpuid240])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc240_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid240/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 240 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid240]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc240_phy_pc_w))
                begin
                    if(good[long_cpuid240/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid240 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid240/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid240])
        end // if (done[240])

        if (done[241]) begin
            timeout[long_cpuid241] = 0;
            //check_bad_trap(spc241_phy_pc_w, 241, long_cpuid241);
            if(active_thread[long_cpuid241])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc241_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid241/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 241 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid241]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc241_phy_pc_w))
                begin
                    if(good[long_cpuid241/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid241 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid241/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid241])
        end // if (done[241])

        if (done[242]) begin
            timeout[long_cpuid242] = 0;
            //check_bad_trap(spc242_phy_pc_w, 242, long_cpuid242);
            if(active_thread[long_cpuid242])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc242_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid242/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 242 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid242]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc242_phy_pc_w))
                begin
                    if(good[long_cpuid242/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid242 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid242/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid242])
        end // if (done[242])

        if (done[243]) begin
            timeout[long_cpuid243] = 0;
            //check_bad_trap(spc243_phy_pc_w, 243, long_cpuid243);
            if(active_thread[long_cpuid243])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc243_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid243/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 243 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid243]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc243_phy_pc_w))
                begin
                    if(good[long_cpuid243/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid243 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid243/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid243])
        end // if (done[243])

        if (done[244]) begin
            timeout[long_cpuid244] = 0;
            //check_bad_trap(spc244_phy_pc_w, 244, long_cpuid244);
            if(active_thread[long_cpuid244])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc244_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid244/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 244 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid244]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc244_phy_pc_w))
                begin
                    if(good[long_cpuid244/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid244 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid244/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid244])
        end // if (done[244])

        if (done[245]) begin
            timeout[long_cpuid245] = 0;
            //check_bad_trap(spc245_phy_pc_w, 245, long_cpuid245);
            if(active_thread[long_cpuid245])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc245_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid245/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 245 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid245]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc245_phy_pc_w))
                begin
                    if(good[long_cpuid245/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid245 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid245/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid245])
        end // if (done[245])

        if (done[246]) begin
            timeout[long_cpuid246] = 0;
            //check_bad_trap(spc246_phy_pc_w, 246, long_cpuid246);
            if(active_thread[long_cpuid246])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc246_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid246/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 246 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid246]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc246_phy_pc_w))
                begin
                    if(good[long_cpuid246/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid246 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid246/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid246])
        end // if (done[246])

        if (done[247]) begin
            timeout[long_cpuid247] = 0;
            //check_bad_trap(spc247_phy_pc_w, 247, long_cpuid247);
            if(active_thread[long_cpuid247])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc247_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid247/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 247 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid247]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc247_phy_pc_w))
                begin
                    if(good[long_cpuid247/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid247 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid247/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid247])
        end // if (done[247])

        if (done[248]) begin
            timeout[long_cpuid248] = 0;
            //check_bad_trap(spc248_phy_pc_w, 248, long_cpuid248);
            if(active_thread[long_cpuid248])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc248_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid248/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 248 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid248]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc248_phy_pc_w))
                begin
                    if(good[long_cpuid248/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid248 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid248/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid248])
        end // if (done[248])

        if (done[249]) begin
            timeout[long_cpuid249] = 0;
            //check_bad_trap(spc249_phy_pc_w, 249, long_cpuid249);
            if(active_thread[long_cpuid249])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc249_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid249/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 249 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid249]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc249_phy_pc_w))
                begin
                    if(good[long_cpuid249/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid249 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid249/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid249])
        end // if (done[249])

        if (done[250]) begin
            timeout[long_cpuid250] = 0;
            //check_bad_trap(spc250_phy_pc_w, 250, long_cpuid250);
            if(active_thread[long_cpuid250])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc250_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid250/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 250 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid250]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc250_phy_pc_w))
                begin
                    if(good[long_cpuid250/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid250 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid250/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid250])
        end // if (done[250])

        if (done[251]) begin
            timeout[long_cpuid251] = 0;
            //check_bad_trap(spc251_phy_pc_w, 251, long_cpuid251);
            if(active_thread[long_cpuid251])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc251_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid251/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 251 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid251]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc251_phy_pc_w))
                begin
                    if(good[long_cpuid251/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid251 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid251/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid251])
        end // if (done[251])

        if (done[252]) begin
            timeout[long_cpuid252] = 0;
            //check_bad_trap(spc252_phy_pc_w, 252, long_cpuid252);
            if(active_thread[long_cpuid252])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc252_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid252/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 252 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid252]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc252_phy_pc_w))
                begin
                    if(good[long_cpuid252/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid252 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid252/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid252])
        end // if (done[252])

        if (done[253]) begin
            timeout[long_cpuid253] = 0;
            //check_bad_trap(spc253_phy_pc_w, 253, long_cpuid253);
            if(active_thread[long_cpuid253])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc253_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid253/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 253 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid253]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc253_phy_pc_w))
                begin
                    if(good[long_cpuid253/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid253 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid253/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid253])
        end // if (done[253])

        if (done[254]) begin
            timeout[long_cpuid254] = 0;
            //check_bad_trap(spc254_phy_pc_w, 254, long_cpuid254);
            if(active_thread[long_cpuid254])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc254_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid254/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 254 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid254]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc254_phy_pc_w))
                begin
                    if(good[long_cpuid254/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid254 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid254/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid254])
        end // if (done[254])

        if (done[255]) begin
            timeout[long_cpuid255] = 0;
            //check_bad_trap(spc255_phy_pc_w, 255, long_cpuid255);
            if(active_thread[long_cpuid255])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc255_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid255/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 255 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid255]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc255_phy_pc_w))
                begin
                    if(good[long_cpuid255/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid255 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid255/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid255])
        end // if (done[255])

        if (done[256]) begin
            timeout[long_cpuid256] = 0;
            //check_bad_trap(spc256_phy_pc_w, 256, long_cpuid256);
            if(active_thread[long_cpuid256])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc256_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid256/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 256 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid256]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc256_phy_pc_w))
                begin
                    if(good[long_cpuid256/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid256 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid256/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid256])
        end // if (done[256])

        if (done[257]) begin
            timeout[long_cpuid257] = 0;
            //check_bad_trap(spc257_phy_pc_w, 257, long_cpuid257);
            if(active_thread[long_cpuid257])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc257_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid257/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 257 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid257]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc257_phy_pc_w))
                begin
                    if(good[long_cpuid257/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid257 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid257/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid257])
        end // if (done[257])

        if (done[258]) begin
            timeout[long_cpuid258] = 0;
            //check_bad_trap(spc258_phy_pc_w, 258, long_cpuid258);
            if(active_thread[long_cpuid258])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc258_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid258/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 258 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid258]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc258_phy_pc_w))
                begin
                    if(good[long_cpuid258/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid258 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid258/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid258])
        end // if (done[258])

        if (done[259]) begin
            timeout[long_cpuid259] = 0;
            //check_bad_trap(spc259_phy_pc_w, 259, long_cpuid259);
            if(active_thread[long_cpuid259])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc259_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid259/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 259 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid259]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc259_phy_pc_w))
                begin
                    if(good[long_cpuid259/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid259 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid259/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid259])
        end // if (done[259])

        if (done[260]) begin
            timeout[long_cpuid260] = 0;
            //check_bad_trap(spc260_phy_pc_w, 260, long_cpuid260);
            if(active_thread[long_cpuid260])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc260_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid260/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 260 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid260]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc260_phy_pc_w))
                begin
                    if(good[long_cpuid260/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid260 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid260/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid260])
        end // if (done[260])

        if (done[261]) begin
            timeout[long_cpuid261] = 0;
            //check_bad_trap(spc261_phy_pc_w, 261, long_cpuid261);
            if(active_thread[long_cpuid261])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc261_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid261/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 261 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid261]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc261_phy_pc_w))
                begin
                    if(good[long_cpuid261/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid261 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid261/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid261])
        end // if (done[261])

        if (done[262]) begin
            timeout[long_cpuid262] = 0;
            //check_bad_trap(spc262_phy_pc_w, 262, long_cpuid262);
            if(active_thread[long_cpuid262])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc262_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid262/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 262 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid262]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc262_phy_pc_w))
                begin
                    if(good[long_cpuid262/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid262 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid262/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid262])
        end // if (done[262])

        if (done[263]) begin
            timeout[long_cpuid263] = 0;
            //check_bad_trap(spc263_phy_pc_w, 263, long_cpuid263);
            if(active_thread[long_cpuid263])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc263_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid263/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 263 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid263]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc263_phy_pc_w))
                begin
                    if(good[long_cpuid263/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid263 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid263/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid263])
        end // if (done[263])

        if (done[264]) begin
            timeout[long_cpuid264] = 0;
            //check_bad_trap(spc264_phy_pc_w, 264, long_cpuid264);
            if(active_thread[long_cpuid264])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc264_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid264/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 264 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid264]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc264_phy_pc_w))
                begin
                    if(good[long_cpuid264/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid264 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid264/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid264])
        end // if (done[264])

        if (done[265]) begin
            timeout[long_cpuid265] = 0;
            //check_bad_trap(spc265_phy_pc_w, 265, long_cpuid265);
            if(active_thread[long_cpuid265])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc265_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid265/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 265 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid265]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc265_phy_pc_w))
                begin
                    if(good[long_cpuid265/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid265 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid265/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid265])
        end // if (done[265])

        if (done[266]) begin
            timeout[long_cpuid266] = 0;
            //check_bad_trap(spc266_phy_pc_w, 266, long_cpuid266);
            if(active_thread[long_cpuid266])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc266_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid266/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 266 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid266]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc266_phy_pc_w))
                begin
                    if(good[long_cpuid266/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid266 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid266/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid266])
        end // if (done[266])

        if (done[267]) begin
            timeout[long_cpuid267] = 0;
            //check_bad_trap(spc267_phy_pc_w, 267, long_cpuid267);
            if(active_thread[long_cpuid267])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc267_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid267/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 267 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid267]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc267_phy_pc_w))
                begin
                    if(good[long_cpuid267/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid267 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid267/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid267])
        end // if (done[267])

        if (done[268]) begin
            timeout[long_cpuid268] = 0;
            //check_bad_trap(spc268_phy_pc_w, 268, long_cpuid268);
            if(active_thread[long_cpuid268])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc268_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid268/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 268 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid268]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc268_phy_pc_w))
                begin
                    if(good[long_cpuid268/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid268 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid268/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid268])
        end // if (done[268])

        if (done[269]) begin
            timeout[long_cpuid269] = 0;
            //check_bad_trap(spc269_phy_pc_w, 269, long_cpuid269);
            if(active_thread[long_cpuid269])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc269_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid269/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 269 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid269]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc269_phy_pc_w))
                begin
                    if(good[long_cpuid269/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid269 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid269/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid269])
        end // if (done[269])

        if (done[270]) begin
            timeout[long_cpuid270] = 0;
            //check_bad_trap(spc270_phy_pc_w, 270, long_cpuid270);
            if(active_thread[long_cpuid270])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc270_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid270/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 270 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid270]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc270_phy_pc_w))
                begin
                    if(good[long_cpuid270/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid270 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid270/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid270])
        end // if (done[270])

        if (done[271]) begin
            timeout[long_cpuid271] = 0;
            //check_bad_trap(spc271_phy_pc_w, 271, long_cpuid271);
            if(active_thread[long_cpuid271])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc271_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid271/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 271 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid271]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc271_phy_pc_w))
                begin
                    if(good[long_cpuid271/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid271 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid271/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid271])
        end // if (done[271])

        if (done[272]) begin
            timeout[long_cpuid272] = 0;
            //check_bad_trap(spc272_phy_pc_w, 272, long_cpuid272);
            if(active_thread[long_cpuid272])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc272_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid272/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 272 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid272]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc272_phy_pc_w))
                begin
                    if(good[long_cpuid272/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid272 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid272/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid272])
        end // if (done[272])

        if (done[273]) begin
            timeout[long_cpuid273] = 0;
            //check_bad_trap(spc273_phy_pc_w, 273, long_cpuid273);
            if(active_thread[long_cpuid273])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc273_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid273/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 273 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid273]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc273_phy_pc_w))
                begin
                    if(good[long_cpuid273/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid273 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid273/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid273])
        end // if (done[273])

        if (done[274]) begin
            timeout[long_cpuid274] = 0;
            //check_bad_trap(spc274_phy_pc_w, 274, long_cpuid274);
            if(active_thread[long_cpuid274])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc274_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid274/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 274 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid274]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc274_phy_pc_w))
                begin
                    if(good[long_cpuid274/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid274 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid274/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid274])
        end // if (done[274])

        if (done[275]) begin
            timeout[long_cpuid275] = 0;
            //check_bad_trap(spc275_phy_pc_w, 275, long_cpuid275);
            if(active_thread[long_cpuid275])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc275_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid275/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 275 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid275]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc275_phy_pc_w))
                begin
                    if(good[long_cpuid275/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid275 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid275/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid275])
        end // if (done[275])

        if (done[276]) begin
            timeout[long_cpuid276] = 0;
            //check_bad_trap(spc276_phy_pc_w, 276, long_cpuid276);
            if(active_thread[long_cpuid276])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc276_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid276/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 276 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid276]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc276_phy_pc_w))
                begin
                    if(good[long_cpuid276/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid276 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid276/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid276])
        end // if (done[276])

        if (done[277]) begin
            timeout[long_cpuid277] = 0;
            //check_bad_trap(spc277_phy_pc_w, 277, long_cpuid277);
            if(active_thread[long_cpuid277])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc277_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid277/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 277 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid277]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc277_phy_pc_w))
                begin
                    if(good[long_cpuid277/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid277 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid277/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid277])
        end // if (done[277])

        if (done[278]) begin
            timeout[long_cpuid278] = 0;
            //check_bad_trap(spc278_phy_pc_w, 278, long_cpuid278);
            if(active_thread[long_cpuid278])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc278_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid278/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 278 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid278]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc278_phy_pc_w))
                begin
                    if(good[long_cpuid278/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid278 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid278/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid278])
        end // if (done[278])

        if (done[279]) begin
            timeout[long_cpuid279] = 0;
            //check_bad_trap(spc279_phy_pc_w, 279, long_cpuid279);
            if(active_thread[long_cpuid279])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc279_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid279/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 279 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid279]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc279_phy_pc_w))
                begin
                    if(good[long_cpuid279/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid279 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid279/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid279])
        end // if (done[279])

        if (done[280]) begin
            timeout[long_cpuid280] = 0;
            //check_bad_trap(spc280_phy_pc_w, 280, long_cpuid280);
            if(active_thread[long_cpuid280])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc280_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid280/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 280 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid280]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc280_phy_pc_w))
                begin
                    if(good[long_cpuid280/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid280 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid280/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid280])
        end // if (done[280])

        if (done[281]) begin
            timeout[long_cpuid281] = 0;
            //check_bad_trap(spc281_phy_pc_w, 281, long_cpuid281);
            if(active_thread[long_cpuid281])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc281_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid281/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 281 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid281]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc281_phy_pc_w))
                begin
                    if(good[long_cpuid281/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid281 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid281/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid281])
        end // if (done[281])

        if (done[282]) begin
            timeout[long_cpuid282] = 0;
            //check_bad_trap(spc282_phy_pc_w, 282, long_cpuid282);
            if(active_thread[long_cpuid282])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc282_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid282/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 282 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid282]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc282_phy_pc_w))
                begin
                    if(good[long_cpuid282/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid282 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid282/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid282])
        end // if (done[282])

        if (done[283]) begin
            timeout[long_cpuid283] = 0;
            //check_bad_trap(spc283_phy_pc_w, 283, long_cpuid283);
            if(active_thread[long_cpuid283])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc283_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid283/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 283 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid283]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc283_phy_pc_w))
                begin
                    if(good[long_cpuid283/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid283 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid283/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid283])
        end // if (done[283])

        if (done[284]) begin
            timeout[long_cpuid284] = 0;
            //check_bad_trap(spc284_phy_pc_w, 284, long_cpuid284);
            if(active_thread[long_cpuid284])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc284_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid284/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 284 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid284]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc284_phy_pc_w))
                begin
                    if(good[long_cpuid284/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid284 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid284/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid284])
        end // if (done[284])

        if (done[285]) begin
            timeout[long_cpuid285] = 0;
            //check_bad_trap(spc285_phy_pc_w, 285, long_cpuid285);
            if(active_thread[long_cpuid285])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc285_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid285/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 285 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid285]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc285_phy_pc_w))
                begin
                    if(good[long_cpuid285/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid285 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid285/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid285])
        end // if (done[285])

        if (done[286]) begin
            timeout[long_cpuid286] = 0;
            //check_bad_trap(spc286_phy_pc_w, 286, long_cpuid286);
            if(active_thread[long_cpuid286])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc286_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid286/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 286 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid286]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc286_phy_pc_w))
                begin
                    if(good[long_cpuid286/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid286 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid286/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid286])
        end // if (done[286])

        if (done[287]) begin
            timeout[long_cpuid287] = 0;
            //check_bad_trap(spc287_phy_pc_w, 287, long_cpuid287);
            if(active_thread[long_cpuid287])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc287_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid287/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 287 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid287]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc287_phy_pc_w))
                begin
                    if(good[long_cpuid287/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid287 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid287/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid287])
        end // if (done[287])

        if (done[288]) begin
            timeout[long_cpuid288] = 0;
            //check_bad_trap(spc288_phy_pc_w, 288, long_cpuid288);
            if(active_thread[long_cpuid288])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc288_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid288/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 288 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid288]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc288_phy_pc_w))
                begin
                    if(good[long_cpuid288/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid288 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid288/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid288])
        end // if (done[288])

        if (done[289]) begin
            timeout[long_cpuid289] = 0;
            //check_bad_trap(spc289_phy_pc_w, 289, long_cpuid289);
            if(active_thread[long_cpuid289])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc289_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid289/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 289 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid289]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc289_phy_pc_w))
                begin
                    if(good[long_cpuid289/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid289 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid289/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid289])
        end // if (done[289])

        if (done[290]) begin
            timeout[long_cpuid290] = 0;
            //check_bad_trap(spc290_phy_pc_w, 290, long_cpuid290);
            if(active_thread[long_cpuid290])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc290_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid290/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 290 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid290]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc290_phy_pc_w))
                begin
                    if(good[long_cpuid290/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid290 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid290/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid290])
        end // if (done[290])

        if (done[291]) begin
            timeout[long_cpuid291] = 0;
            //check_bad_trap(spc291_phy_pc_w, 291, long_cpuid291);
            if(active_thread[long_cpuid291])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc291_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid291/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 291 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid291]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc291_phy_pc_w))
                begin
                    if(good[long_cpuid291/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid291 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid291/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid291])
        end // if (done[291])

        if (done[292]) begin
            timeout[long_cpuid292] = 0;
            //check_bad_trap(spc292_phy_pc_w, 292, long_cpuid292);
            if(active_thread[long_cpuid292])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc292_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid292/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 292 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid292]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc292_phy_pc_w))
                begin
                    if(good[long_cpuid292/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid292 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid292/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid292])
        end // if (done[292])

        if (done[293]) begin
            timeout[long_cpuid293] = 0;
            //check_bad_trap(spc293_phy_pc_w, 293, long_cpuid293);
            if(active_thread[long_cpuid293])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc293_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid293/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 293 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid293]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc293_phy_pc_w))
                begin
                    if(good[long_cpuid293/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid293 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid293/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid293])
        end // if (done[293])

        if (done[294]) begin
            timeout[long_cpuid294] = 0;
            //check_bad_trap(spc294_phy_pc_w, 294, long_cpuid294);
            if(active_thread[long_cpuid294])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc294_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid294/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 294 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid294]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc294_phy_pc_w))
                begin
                    if(good[long_cpuid294/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid294 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid294/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid294])
        end // if (done[294])

        if (done[295]) begin
            timeout[long_cpuid295] = 0;
            //check_bad_trap(spc295_phy_pc_w, 295, long_cpuid295);
            if(active_thread[long_cpuid295])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc295_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid295/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 295 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid295]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc295_phy_pc_w))
                begin
                    if(good[long_cpuid295/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid295 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid295/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid295])
        end // if (done[295])

        if (done[296]) begin
            timeout[long_cpuid296] = 0;
            //check_bad_trap(spc296_phy_pc_w, 296, long_cpuid296);
            if(active_thread[long_cpuid296])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc296_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid296/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 296 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid296]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc296_phy_pc_w))
                begin
                    if(good[long_cpuid296/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid296 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid296/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid296])
        end // if (done[296])

        if (done[297]) begin
            timeout[long_cpuid297] = 0;
            //check_bad_trap(spc297_phy_pc_w, 297, long_cpuid297);
            if(active_thread[long_cpuid297])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc297_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid297/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 297 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid297]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc297_phy_pc_w))
                begin
                    if(good[long_cpuid297/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid297 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid297/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid297])
        end // if (done[297])

        if (done[298]) begin
            timeout[long_cpuid298] = 0;
            //check_bad_trap(spc298_phy_pc_w, 298, long_cpuid298);
            if(active_thread[long_cpuid298])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc298_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid298/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 298 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid298]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc298_phy_pc_w))
                begin
                    if(good[long_cpuid298/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid298 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid298/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid298])
        end // if (done[298])

        if (done[299]) begin
            timeout[long_cpuid299] = 0;
            //check_bad_trap(spc299_phy_pc_w, 299, long_cpuid299);
            if(active_thread[long_cpuid299])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc299_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid299/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 299 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid299]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc299_phy_pc_w))
                begin
                    if(good[long_cpuid299/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid299 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid299/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid299])
        end // if (done[299])

        if (done[300]) begin
            timeout[long_cpuid300] = 0;
            //check_bad_trap(spc300_phy_pc_w, 300, long_cpuid300);
            if(active_thread[long_cpuid300])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc300_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid300/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 300 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid300]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc300_phy_pc_w))
                begin
                    if(good[long_cpuid300/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid300 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid300/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid300])
        end // if (done[300])

        if (done[301]) begin
            timeout[long_cpuid301] = 0;
            //check_bad_trap(spc301_phy_pc_w, 301, long_cpuid301);
            if(active_thread[long_cpuid301])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc301_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid301/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 301 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid301]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc301_phy_pc_w))
                begin
                    if(good[long_cpuid301/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid301 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid301/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid301])
        end // if (done[301])

        if (done[302]) begin
            timeout[long_cpuid302] = 0;
            //check_bad_trap(spc302_phy_pc_w, 302, long_cpuid302);
            if(active_thread[long_cpuid302])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc302_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid302/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 302 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid302]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc302_phy_pc_w))
                begin
                    if(good[long_cpuid302/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid302 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid302/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid302])
        end // if (done[302])

        if (done[303]) begin
            timeout[long_cpuid303] = 0;
            //check_bad_trap(spc303_phy_pc_w, 303, long_cpuid303);
            if(active_thread[long_cpuid303])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc303_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid303/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 303 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid303]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc303_phy_pc_w))
                begin
                    if(good[long_cpuid303/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid303 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid303/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid303])
        end // if (done[303])

        if (done[304]) begin
            timeout[long_cpuid304] = 0;
            //check_bad_trap(spc304_phy_pc_w, 304, long_cpuid304);
            if(active_thread[long_cpuid304])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc304_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid304/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 304 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid304]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc304_phy_pc_w))
                begin
                    if(good[long_cpuid304/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid304 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid304/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid304])
        end // if (done[304])

        if (done[305]) begin
            timeout[long_cpuid305] = 0;
            //check_bad_trap(spc305_phy_pc_w, 305, long_cpuid305);
            if(active_thread[long_cpuid305])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc305_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid305/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 305 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid305]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc305_phy_pc_w))
                begin
                    if(good[long_cpuid305/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid305 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid305/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid305])
        end // if (done[305])

        if (done[306]) begin
            timeout[long_cpuid306] = 0;
            //check_bad_trap(spc306_phy_pc_w, 306, long_cpuid306);
            if(active_thread[long_cpuid306])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc306_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid306/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 306 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid306]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc306_phy_pc_w))
                begin
                    if(good[long_cpuid306/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid306 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid306/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid306])
        end // if (done[306])

        if (done[307]) begin
            timeout[long_cpuid307] = 0;
            //check_bad_trap(spc307_phy_pc_w, 307, long_cpuid307);
            if(active_thread[long_cpuid307])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc307_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid307/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 307 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid307]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc307_phy_pc_w))
                begin
                    if(good[long_cpuid307/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid307 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid307/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid307])
        end // if (done[307])

        if (done[308]) begin
            timeout[long_cpuid308] = 0;
            //check_bad_trap(spc308_phy_pc_w, 308, long_cpuid308);
            if(active_thread[long_cpuid308])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc308_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid308/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 308 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid308]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc308_phy_pc_w))
                begin
                    if(good[long_cpuid308/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid308 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid308/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid308])
        end // if (done[308])

        if (done[309]) begin
            timeout[long_cpuid309] = 0;
            //check_bad_trap(spc309_phy_pc_w, 309, long_cpuid309);
            if(active_thread[long_cpuid309])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc309_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid309/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 309 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid309]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc309_phy_pc_w))
                begin
                    if(good[long_cpuid309/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid309 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid309/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid309])
        end // if (done[309])

        if (done[310]) begin
            timeout[long_cpuid310] = 0;
            //check_bad_trap(spc310_phy_pc_w, 310, long_cpuid310);
            if(active_thread[long_cpuid310])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc310_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid310/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 310 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid310]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc310_phy_pc_w))
                begin
                    if(good[long_cpuid310/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid310 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid310/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid310])
        end // if (done[310])

        if (done[311]) begin
            timeout[long_cpuid311] = 0;
            //check_bad_trap(spc311_phy_pc_w, 311, long_cpuid311);
            if(active_thread[long_cpuid311])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc311_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid311/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 311 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid311]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc311_phy_pc_w))
                begin
                    if(good[long_cpuid311/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid311 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid311/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid311])
        end // if (done[311])

        if (done[312]) begin
            timeout[long_cpuid312] = 0;
            //check_bad_trap(spc312_phy_pc_w, 312, long_cpuid312);
            if(active_thread[long_cpuid312])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc312_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid312/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 312 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid312]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc312_phy_pc_w))
                begin
                    if(good[long_cpuid312/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid312 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid312/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid312])
        end // if (done[312])

        if (done[313]) begin
            timeout[long_cpuid313] = 0;
            //check_bad_trap(spc313_phy_pc_w, 313, long_cpuid313);
            if(active_thread[long_cpuid313])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc313_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid313/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 313 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid313]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc313_phy_pc_w))
                begin
                    if(good[long_cpuid313/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid313 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid313/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid313])
        end // if (done[313])

        if (done[314]) begin
            timeout[long_cpuid314] = 0;
            //check_bad_trap(spc314_phy_pc_w, 314, long_cpuid314);
            if(active_thread[long_cpuid314])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc314_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid314/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 314 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid314]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc314_phy_pc_w))
                begin
                    if(good[long_cpuid314/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid314 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid314/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid314])
        end // if (done[314])

        if (done[315]) begin
            timeout[long_cpuid315] = 0;
            //check_bad_trap(spc315_phy_pc_w, 315, long_cpuid315);
            if(active_thread[long_cpuid315])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc315_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid315/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 315 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid315]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc315_phy_pc_w))
                begin
                    if(good[long_cpuid315/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid315 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid315/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid315])
        end // if (done[315])

        if (done[316]) begin
            timeout[long_cpuid316] = 0;
            //check_bad_trap(spc316_phy_pc_w, 316, long_cpuid316);
            if(active_thread[long_cpuid316])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc316_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid316/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 316 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid316]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc316_phy_pc_w))
                begin
                    if(good[long_cpuid316/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid316 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid316/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid316])
        end // if (done[316])

        if (done[317]) begin
            timeout[long_cpuid317] = 0;
            //check_bad_trap(spc317_phy_pc_w, 317, long_cpuid317);
            if(active_thread[long_cpuid317])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc317_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid317/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 317 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid317]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc317_phy_pc_w))
                begin
                    if(good[long_cpuid317/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid317 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid317/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid317])
        end // if (done[317])

        if (done[318]) begin
            timeout[long_cpuid318] = 0;
            //check_bad_trap(spc318_phy_pc_w, 318, long_cpuid318);
            if(active_thread[long_cpuid318])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc318_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid318/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 318 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid318]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc318_phy_pc_w))
                begin
                    if(good[long_cpuid318/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid318 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid318/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid318])
        end // if (done[318])

        if (done[319]) begin
            timeout[long_cpuid319] = 0;
            //check_bad_trap(spc319_phy_pc_w, 319, long_cpuid319);
            if(active_thread[long_cpuid319])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc319_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid319/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 319 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid319]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc319_phy_pc_w))
                begin
                    if(good[long_cpuid319/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid319 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid319/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid319])
        end // if (done[319])

        if (done[320]) begin
            timeout[long_cpuid320] = 0;
            //check_bad_trap(spc320_phy_pc_w, 320, long_cpuid320);
            if(active_thread[long_cpuid320])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc320_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid320/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 320 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid320]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc320_phy_pc_w))
                begin
                    if(good[long_cpuid320/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid320 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid320/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid320])
        end // if (done[320])

        if (done[321]) begin
            timeout[long_cpuid321] = 0;
            //check_bad_trap(spc321_phy_pc_w, 321, long_cpuid321);
            if(active_thread[long_cpuid321])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc321_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid321/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 321 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid321]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc321_phy_pc_w))
                begin
                    if(good[long_cpuid321/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid321 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid321/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid321])
        end // if (done[321])

        if (done[322]) begin
            timeout[long_cpuid322] = 0;
            //check_bad_trap(spc322_phy_pc_w, 322, long_cpuid322);
            if(active_thread[long_cpuid322])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc322_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid322/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 322 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid322]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc322_phy_pc_w))
                begin
                    if(good[long_cpuid322/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid322 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid322/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid322])
        end // if (done[322])

        if (done[323]) begin
            timeout[long_cpuid323] = 0;
            //check_bad_trap(spc323_phy_pc_w, 323, long_cpuid323);
            if(active_thread[long_cpuid323])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc323_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid323/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 323 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid323]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc323_phy_pc_w))
                begin
                    if(good[long_cpuid323/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid323 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid323/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid323])
        end // if (done[323])

        if (done[324]) begin
            timeout[long_cpuid324] = 0;
            //check_bad_trap(spc324_phy_pc_w, 324, long_cpuid324);
            if(active_thread[long_cpuid324])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc324_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid324/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 324 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid324]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc324_phy_pc_w))
                begin
                    if(good[long_cpuid324/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid324 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid324/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid324])
        end // if (done[324])

        if (done[325]) begin
            timeout[long_cpuid325] = 0;
            //check_bad_trap(spc325_phy_pc_w, 325, long_cpuid325);
            if(active_thread[long_cpuid325])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc325_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid325/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 325 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid325]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc325_phy_pc_w))
                begin
                    if(good[long_cpuid325/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid325 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid325/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid325])
        end // if (done[325])

        if (done[326]) begin
            timeout[long_cpuid326] = 0;
            //check_bad_trap(spc326_phy_pc_w, 326, long_cpuid326);
            if(active_thread[long_cpuid326])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc326_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid326/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 326 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid326]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc326_phy_pc_w))
                begin
                    if(good[long_cpuid326/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid326 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid326/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid326])
        end // if (done[326])

        if (done[327]) begin
            timeout[long_cpuid327] = 0;
            //check_bad_trap(spc327_phy_pc_w, 327, long_cpuid327);
            if(active_thread[long_cpuid327])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc327_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid327/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 327 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid327]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc327_phy_pc_w))
                begin
                    if(good[long_cpuid327/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid327 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid327/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid327])
        end // if (done[327])

        if (done[328]) begin
            timeout[long_cpuid328] = 0;
            //check_bad_trap(spc328_phy_pc_w, 328, long_cpuid328);
            if(active_thread[long_cpuid328])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc328_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid328/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 328 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid328]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc328_phy_pc_w))
                begin
                    if(good[long_cpuid328/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid328 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid328/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid328])
        end // if (done[328])

        if (done[329]) begin
            timeout[long_cpuid329] = 0;
            //check_bad_trap(spc329_phy_pc_w, 329, long_cpuid329);
            if(active_thread[long_cpuid329])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc329_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid329/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 329 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid329]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc329_phy_pc_w))
                begin
                    if(good[long_cpuid329/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid329 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid329/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid329])
        end // if (done[329])

        if (done[330]) begin
            timeout[long_cpuid330] = 0;
            //check_bad_trap(spc330_phy_pc_w, 330, long_cpuid330);
            if(active_thread[long_cpuid330])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc330_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid330/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 330 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid330]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc330_phy_pc_w))
                begin
                    if(good[long_cpuid330/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid330 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid330/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid330])
        end // if (done[330])

        if (done[331]) begin
            timeout[long_cpuid331] = 0;
            //check_bad_trap(spc331_phy_pc_w, 331, long_cpuid331);
            if(active_thread[long_cpuid331])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc331_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid331/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 331 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid331]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc331_phy_pc_w))
                begin
                    if(good[long_cpuid331/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid331 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid331/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid331])
        end // if (done[331])

        if (done[332]) begin
            timeout[long_cpuid332] = 0;
            //check_bad_trap(spc332_phy_pc_w, 332, long_cpuid332);
            if(active_thread[long_cpuid332])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc332_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid332/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 332 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid332]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc332_phy_pc_w))
                begin
                    if(good[long_cpuid332/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid332 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid332/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid332])
        end // if (done[332])

        if (done[333]) begin
            timeout[long_cpuid333] = 0;
            //check_bad_trap(spc333_phy_pc_w, 333, long_cpuid333);
            if(active_thread[long_cpuid333])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc333_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid333/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 333 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid333]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc333_phy_pc_w))
                begin
                    if(good[long_cpuid333/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid333 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid333/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid333])
        end // if (done[333])

        if (done[334]) begin
            timeout[long_cpuid334] = 0;
            //check_bad_trap(spc334_phy_pc_w, 334, long_cpuid334);
            if(active_thread[long_cpuid334])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc334_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid334/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 334 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid334]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc334_phy_pc_w))
                begin
                    if(good[long_cpuid334/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid334 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid334/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid334])
        end // if (done[334])

        if (done[335]) begin
            timeout[long_cpuid335] = 0;
            //check_bad_trap(spc335_phy_pc_w, 335, long_cpuid335);
            if(active_thread[long_cpuid335])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc335_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid335/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 335 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid335]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc335_phy_pc_w))
                begin
                    if(good[long_cpuid335/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid335 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid335/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid335])
        end // if (done[335])

        if (done[336]) begin
            timeout[long_cpuid336] = 0;
            //check_bad_trap(spc336_phy_pc_w, 336, long_cpuid336);
            if(active_thread[long_cpuid336])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc336_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid336/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 336 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid336]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc336_phy_pc_w))
                begin
                    if(good[long_cpuid336/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid336 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid336/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid336])
        end // if (done[336])

        if (done[337]) begin
            timeout[long_cpuid337] = 0;
            //check_bad_trap(spc337_phy_pc_w, 337, long_cpuid337);
            if(active_thread[long_cpuid337])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc337_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid337/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 337 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid337]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc337_phy_pc_w))
                begin
                    if(good[long_cpuid337/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid337 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid337/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid337])
        end // if (done[337])

        if (done[338]) begin
            timeout[long_cpuid338] = 0;
            //check_bad_trap(spc338_phy_pc_w, 338, long_cpuid338);
            if(active_thread[long_cpuid338])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc338_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid338/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 338 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid338]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc338_phy_pc_w))
                begin
                    if(good[long_cpuid338/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid338 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid338/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid338])
        end // if (done[338])

        if (done[339]) begin
            timeout[long_cpuid339] = 0;
            //check_bad_trap(spc339_phy_pc_w, 339, long_cpuid339);
            if(active_thread[long_cpuid339])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc339_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid339/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 339 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid339]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc339_phy_pc_w))
                begin
                    if(good[long_cpuid339/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid339 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid339/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid339])
        end // if (done[339])

        if (done[340]) begin
            timeout[long_cpuid340] = 0;
            //check_bad_trap(spc340_phy_pc_w, 340, long_cpuid340);
            if(active_thread[long_cpuid340])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc340_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid340/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 340 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid340]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc340_phy_pc_w))
                begin
                    if(good[long_cpuid340/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid340 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid340/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid340])
        end // if (done[340])

        if (done[341]) begin
            timeout[long_cpuid341] = 0;
            //check_bad_trap(spc341_phy_pc_w, 341, long_cpuid341);
            if(active_thread[long_cpuid341])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc341_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid341/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 341 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid341]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc341_phy_pc_w))
                begin
                    if(good[long_cpuid341/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid341 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid341/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid341])
        end // if (done[341])

        if (done[342]) begin
            timeout[long_cpuid342] = 0;
            //check_bad_trap(spc342_phy_pc_w, 342, long_cpuid342);
            if(active_thread[long_cpuid342])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc342_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid342/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 342 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid342]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc342_phy_pc_w))
                begin
                    if(good[long_cpuid342/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid342 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid342/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid342])
        end // if (done[342])

        if (done[343]) begin
            timeout[long_cpuid343] = 0;
            //check_bad_trap(spc343_phy_pc_w, 343, long_cpuid343);
            if(active_thread[long_cpuid343])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc343_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid343/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 343 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid343]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc343_phy_pc_w))
                begin
                    if(good[long_cpuid343/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid343 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid343/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid343])
        end // if (done[343])

        if (done[344]) begin
            timeout[long_cpuid344] = 0;
            //check_bad_trap(spc344_phy_pc_w, 344, long_cpuid344);
            if(active_thread[long_cpuid344])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc344_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid344/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 344 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid344]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc344_phy_pc_w))
                begin
                    if(good[long_cpuid344/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid344 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid344/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid344])
        end // if (done[344])

        if (done[345]) begin
            timeout[long_cpuid345] = 0;
            //check_bad_trap(spc345_phy_pc_w, 345, long_cpuid345);
            if(active_thread[long_cpuid345])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc345_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid345/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 345 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid345]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc345_phy_pc_w))
                begin
                    if(good[long_cpuid345/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid345 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid345/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid345])
        end // if (done[345])

        if (done[346]) begin
            timeout[long_cpuid346] = 0;
            //check_bad_trap(spc346_phy_pc_w, 346, long_cpuid346);
            if(active_thread[long_cpuid346])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc346_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid346/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 346 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid346]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc346_phy_pc_w))
                begin
                    if(good[long_cpuid346/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid346 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid346/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid346])
        end // if (done[346])

        if (done[347]) begin
            timeout[long_cpuid347] = 0;
            //check_bad_trap(spc347_phy_pc_w, 347, long_cpuid347);
            if(active_thread[long_cpuid347])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc347_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid347/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 347 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid347]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc347_phy_pc_w))
                begin
                    if(good[long_cpuid347/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid347 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid347/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid347])
        end // if (done[347])

        if (done[348]) begin
            timeout[long_cpuid348] = 0;
            //check_bad_trap(spc348_phy_pc_w, 348, long_cpuid348);
            if(active_thread[long_cpuid348])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc348_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid348/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 348 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid348]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc348_phy_pc_w))
                begin
                    if(good[long_cpuid348/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid348 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid348/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid348])
        end // if (done[348])

        if (done[349]) begin
            timeout[long_cpuid349] = 0;
            //check_bad_trap(spc349_phy_pc_w, 349, long_cpuid349);
            if(active_thread[long_cpuid349])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc349_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid349/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 349 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid349]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc349_phy_pc_w))
                begin
                    if(good[long_cpuid349/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid349 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid349/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid349])
        end // if (done[349])

        if (done[350]) begin
            timeout[long_cpuid350] = 0;
            //check_bad_trap(spc350_phy_pc_w, 350, long_cpuid350);
            if(active_thread[long_cpuid350])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc350_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid350/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 350 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid350]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc350_phy_pc_w))
                begin
                    if(good[long_cpuid350/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid350 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid350/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid350])
        end // if (done[350])

        if (done[351]) begin
            timeout[long_cpuid351] = 0;
            //check_bad_trap(spc351_phy_pc_w, 351, long_cpuid351);
            if(active_thread[long_cpuid351])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc351_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid351/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 351 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid351]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc351_phy_pc_w))
                begin
                    if(good[long_cpuid351/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid351 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid351/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid351])
        end // if (done[351])

        if (done[352]) begin
            timeout[long_cpuid352] = 0;
            //check_bad_trap(spc352_phy_pc_w, 352, long_cpuid352);
            if(active_thread[long_cpuid352])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc352_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid352/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 352 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid352]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc352_phy_pc_w))
                begin
                    if(good[long_cpuid352/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid352 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid352/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid352])
        end // if (done[352])

        if (done[353]) begin
            timeout[long_cpuid353] = 0;
            //check_bad_trap(spc353_phy_pc_w, 353, long_cpuid353);
            if(active_thread[long_cpuid353])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc353_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid353/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 353 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid353]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc353_phy_pc_w))
                begin
                    if(good[long_cpuid353/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid353 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid353/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid353])
        end // if (done[353])

        if (done[354]) begin
            timeout[long_cpuid354] = 0;
            //check_bad_trap(spc354_phy_pc_w, 354, long_cpuid354);
            if(active_thread[long_cpuid354])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc354_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid354/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 354 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid354]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc354_phy_pc_w))
                begin
                    if(good[long_cpuid354/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid354 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid354/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid354])
        end // if (done[354])

        if (done[355]) begin
            timeout[long_cpuid355] = 0;
            //check_bad_trap(spc355_phy_pc_w, 355, long_cpuid355);
            if(active_thread[long_cpuid355])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc355_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid355/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 355 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid355]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc355_phy_pc_w))
                begin
                    if(good[long_cpuid355/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid355 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid355/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid355])
        end // if (done[355])

        if (done[356]) begin
            timeout[long_cpuid356] = 0;
            //check_bad_trap(spc356_phy_pc_w, 356, long_cpuid356);
            if(active_thread[long_cpuid356])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc356_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid356/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 356 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid356]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc356_phy_pc_w))
                begin
                    if(good[long_cpuid356/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid356 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid356/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid356])
        end // if (done[356])

        if (done[357]) begin
            timeout[long_cpuid357] = 0;
            //check_bad_trap(spc357_phy_pc_w, 357, long_cpuid357);
            if(active_thread[long_cpuid357])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc357_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid357/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 357 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid357]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc357_phy_pc_w))
                begin
                    if(good[long_cpuid357/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid357 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid357/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid357])
        end // if (done[357])

        if (done[358]) begin
            timeout[long_cpuid358] = 0;
            //check_bad_trap(spc358_phy_pc_w, 358, long_cpuid358);
            if(active_thread[long_cpuid358])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc358_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid358/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 358 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid358]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc358_phy_pc_w))
                begin
                    if(good[long_cpuid358/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid358 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid358/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid358])
        end // if (done[358])

        if (done[359]) begin
            timeout[long_cpuid359] = 0;
            //check_bad_trap(spc359_phy_pc_w, 359, long_cpuid359);
            if(active_thread[long_cpuid359])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc359_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid359/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 359 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid359]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc359_phy_pc_w))
                begin
                    if(good[long_cpuid359/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid359 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid359/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid359])
        end // if (done[359])

        if (done[360]) begin
            timeout[long_cpuid360] = 0;
            //check_bad_trap(spc360_phy_pc_w, 360, long_cpuid360);
            if(active_thread[long_cpuid360])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc360_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid360/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 360 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid360]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc360_phy_pc_w))
                begin
                    if(good[long_cpuid360/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid360 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid360/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid360])
        end // if (done[360])

        if (done[361]) begin
            timeout[long_cpuid361] = 0;
            //check_bad_trap(spc361_phy_pc_w, 361, long_cpuid361);
            if(active_thread[long_cpuid361])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc361_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid361/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 361 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid361]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc361_phy_pc_w))
                begin
                    if(good[long_cpuid361/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid361 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid361/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid361])
        end // if (done[361])

        if (done[362]) begin
            timeout[long_cpuid362] = 0;
            //check_bad_trap(spc362_phy_pc_w, 362, long_cpuid362);
            if(active_thread[long_cpuid362])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc362_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid362/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 362 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid362]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc362_phy_pc_w))
                begin
                    if(good[long_cpuid362/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid362 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid362/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid362])
        end // if (done[362])

        if (done[363]) begin
            timeout[long_cpuid363] = 0;
            //check_bad_trap(spc363_phy_pc_w, 363, long_cpuid363);
            if(active_thread[long_cpuid363])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc363_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid363/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 363 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid363]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc363_phy_pc_w))
                begin
                    if(good[long_cpuid363/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid363 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid363/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid363])
        end // if (done[363])

        if (done[364]) begin
            timeout[long_cpuid364] = 0;
            //check_bad_trap(spc364_phy_pc_w, 364, long_cpuid364);
            if(active_thread[long_cpuid364])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc364_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid364/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 364 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid364]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc364_phy_pc_w))
                begin
                    if(good[long_cpuid364/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid364 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid364/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid364])
        end // if (done[364])

        if (done[365]) begin
            timeout[long_cpuid365] = 0;
            //check_bad_trap(spc365_phy_pc_w, 365, long_cpuid365);
            if(active_thread[long_cpuid365])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc365_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid365/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 365 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid365]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc365_phy_pc_w))
                begin
                    if(good[long_cpuid365/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid365 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid365/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid365])
        end // if (done[365])

        if (done[366]) begin
            timeout[long_cpuid366] = 0;
            //check_bad_trap(spc366_phy_pc_w, 366, long_cpuid366);
            if(active_thread[long_cpuid366])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc366_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid366/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 366 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid366]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc366_phy_pc_w))
                begin
                    if(good[long_cpuid366/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid366 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid366/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid366])
        end // if (done[366])

        if (done[367]) begin
            timeout[long_cpuid367] = 0;
            //check_bad_trap(spc367_phy_pc_w, 367, long_cpuid367);
            if(active_thread[long_cpuid367])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc367_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid367/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 367 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid367]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc367_phy_pc_w))
                begin
                    if(good[long_cpuid367/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid367 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid367/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid367])
        end // if (done[367])

        if (done[368]) begin
            timeout[long_cpuid368] = 0;
            //check_bad_trap(spc368_phy_pc_w, 368, long_cpuid368);
            if(active_thread[long_cpuid368])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc368_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid368/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 368 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid368]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc368_phy_pc_w))
                begin
                    if(good[long_cpuid368/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid368 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid368/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid368])
        end // if (done[368])

        if (done[369]) begin
            timeout[long_cpuid369] = 0;
            //check_bad_trap(spc369_phy_pc_w, 369, long_cpuid369);
            if(active_thread[long_cpuid369])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc369_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid369/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 369 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid369]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc369_phy_pc_w))
                begin
                    if(good[long_cpuid369/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid369 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid369/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid369])
        end // if (done[369])

        if (done[370]) begin
            timeout[long_cpuid370] = 0;
            //check_bad_trap(spc370_phy_pc_w, 370, long_cpuid370);
            if(active_thread[long_cpuid370])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc370_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid370/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 370 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid370]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc370_phy_pc_w))
                begin
                    if(good[long_cpuid370/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid370 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid370/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid370])
        end // if (done[370])

        if (done[371]) begin
            timeout[long_cpuid371] = 0;
            //check_bad_trap(spc371_phy_pc_w, 371, long_cpuid371);
            if(active_thread[long_cpuid371])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc371_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid371/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 371 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid371]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc371_phy_pc_w))
                begin
                    if(good[long_cpuid371/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid371 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid371/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid371])
        end // if (done[371])

        if (done[372]) begin
            timeout[long_cpuid372] = 0;
            //check_bad_trap(spc372_phy_pc_w, 372, long_cpuid372);
            if(active_thread[long_cpuid372])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc372_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid372/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 372 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid372]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc372_phy_pc_w))
                begin
                    if(good[long_cpuid372/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid372 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid372/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid372])
        end // if (done[372])

        if (done[373]) begin
            timeout[long_cpuid373] = 0;
            //check_bad_trap(spc373_phy_pc_w, 373, long_cpuid373);
            if(active_thread[long_cpuid373])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc373_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid373/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 373 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid373]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc373_phy_pc_w))
                begin
                    if(good[long_cpuid373/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid373 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid373/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid373])
        end // if (done[373])

        if (done[374]) begin
            timeout[long_cpuid374] = 0;
            //check_bad_trap(spc374_phy_pc_w, 374, long_cpuid374);
            if(active_thread[long_cpuid374])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc374_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid374/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 374 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid374]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc374_phy_pc_w))
                begin
                    if(good[long_cpuid374/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid374 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid374/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid374])
        end // if (done[374])

        if (done[375]) begin
            timeout[long_cpuid375] = 0;
            //check_bad_trap(spc375_phy_pc_w, 375, long_cpuid375);
            if(active_thread[long_cpuid375])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc375_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid375/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 375 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid375]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc375_phy_pc_w))
                begin
                    if(good[long_cpuid375/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid375 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid375/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid375])
        end // if (done[375])

        if (done[376]) begin
            timeout[long_cpuid376] = 0;
            //check_bad_trap(spc376_phy_pc_w, 376, long_cpuid376);
            if(active_thread[long_cpuid376])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc376_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid376/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 376 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid376]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc376_phy_pc_w))
                begin
                    if(good[long_cpuid376/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid376 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid376/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid376])
        end // if (done[376])

        if (done[377]) begin
            timeout[long_cpuid377] = 0;
            //check_bad_trap(spc377_phy_pc_w, 377, long_cpuid377);
            if(active_thread[long_cpuid377])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc377_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid377/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 377 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid377]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc377_phy_pc_w))
                begin
                    if(good[long_cpuid377/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid377 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid377/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid377])
        end // if (done[377])

        if (done[378]) begin
            timeout[long_cpuid378] = 0;
            //check_bad_trap(spc378_phy_pc_w, 378, long_cpuid378);
            if(active_thread[long_cpuid378])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc378_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid378/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 378 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid378]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc378_phy_pc_w))
                begin
                    if(good[long_cpuid378/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid378 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid378/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid378])
        end // if (done[378])

        if (done[379]) begin
            timeout[long_cpuid379] = 0;
            //check_bad_trap(spc379_phy_pc_w, 379, long_cpuid379);
            if(active_thread[long_cpuid379])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc379_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid379/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 379 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid379]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc379_phy_pc_w))
                begin
                    if(good[long_cpuid379/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid379 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid379/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid379])
        end // if (done[379])

        if (done[380]) begin
            timeout[long_cpuid380] = 0;
            //check_bad_trap(spc380_phy_pc_w, 380, long_cpuid380);
            if(active_thread[long_cpuid380])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc380_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid380/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 380 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid380]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc380_phy_pc_w))
                begin
                    if(good[long_cpuid380/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid380 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid380/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid380])
        end // if (done[380])

        if (done[381]) begin
            timeout[long_cpuid381] = 0;
            //check_bad_trap(spc381_phy_pc_w, 381, long_cpuid381);
            if(active_thread[long_cpuid381])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc381_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid381/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 381 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid381]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc381_phy_pc_w))
                begin
                    if(good[long_cpuid381/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid381 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid381/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid381])
        end // if (done[381])

        if (done[382]) begin
            timeout[long_cpuid382] = 0;
            //check_bad_trap(spc382_phy_pc_w, 382, long_cpuid382);
            if(active_thread[long_cpuid382])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc382_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid382/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 382 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid382]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc382_phy_pc_w))
                begin
                    if(good[long_cpuid382/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid382 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid382/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid382])
        end // if (done[382])

        if (done[383]) begin
            timeout[long_cpuid383] = 0;
            //check_bad_trap(spc383_phy_pc_w, 383, long_cpuid383);
            if(active_thread[long_cpuid383])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc383_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid383/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 383 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid383]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc383_phy_pc_w))
                begin
                    if(good[long_cpuid383/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid383 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid383/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid383])
        end // if (done[383])

        if (done[384]) begin
            timeout[long_cpuid384] = 0;
            //check_bad_trap(spc384_phy_pc_w, 384, long_cpuid384);
            if(active_thread[long_cpuid384])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc384_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid384/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 384 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid384]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc384_phy_pc_w))
                begin
                    if(good[long_cpuid384/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid384 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid384/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid384])
        end // if (done[384])

        if (done[385]) begin
            timeout[long_cpuid385] = 0;
            //check_bad_trap(spc385_phy_pc_w, 385, long_cpuid385);
            if(active_thread[long_cpuid385])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc385_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid385/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 385 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid385]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc385_phy_pc_w))
                begin
                    if(good[long_cpuid385/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid385 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid385/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid385])
        end // if (done[385])

        if (done[386]) begin
            timeout[long_cpuid386] = 0;
            //check_bad_trap(spc386_phy_pc_w, 386, long_cpuid386);
            if(active_thread[long_cpuid386])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc386_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid386/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 386 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid386]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc386_phy_pc_w))
                begin
                    if(good[long_cpuid386/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid386 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid386/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid386])
        end // if (done[386])

        if (done[387]) begin
            timeout[long_cpuid387] = 0;
            //check_bad_trap(spc387_phy_pc_w, 387, long_cpuid387);
            if(active_thread[long_cpuid387])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc387_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid387/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 387 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid387]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc387_phy_pc_w))
                begin
                    if(good[long_cpuid387/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid387 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid387/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid387])
        end // if (done[387])

        if (done[388]) begin
            timeout[long_cpuid388] = 0;
            //check_bad_trap(spc388_phy_pc_w, 388, long_cpuid388);
            if(active_thread[long_cpuid388])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc388_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid388/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 388 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid388]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc388_phy_pc_w))
                begin
                    if(good[long_cpuid388/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid388 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid388/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid388])
        end // if (done[388])

        if (done[389]) begin
            timeout[long_cpuid389] = 0;
            //check_bad_trap(spc389_phy_pc_w, 389, long_cpuid389);
            if(active_thread[long_cpuid389])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc389_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid389/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 389 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid389]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc389_phy_pc_w))
                begin
                    if(good[long_cpuid389/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid389 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid389/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid389])
        end // if (done[389])

        if (done[390]) begin
            timeout[long_cpuid390] = 0;
            //check_bad_trap(spc390_phy_pc_w, 390, long_cpuid390);
            if(active_thread[long_cpuid390])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc390_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid390/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 390 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid390]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc390_phy_pc_w))
                begin
                    if(good[long_cpuid390/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid390 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid390/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid390])
        end // if (done[390])

        if (done[391]) begin
            timeout[long_cpuid391] = 0;
            //check_bad_trap(spc391_phy_pc_w, 391, long_cpuid391);
            if(active_thread[long_cpuid391])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc391_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid391/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 391 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid391]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc391_phy_pc_w))
                begin
                    if(good[long_cpuid391/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid391 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid391/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid391])
        end // if (done[391])

        if (done[392]) begin
            timeout[long_cpuid392] = 0;
            //check_bad_trap(spc392_phy_pc_w, 392, long_cpuid392);
            if(active_thread[long_cpuid392])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc392_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid392/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 392 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid392]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc392_phy_pc_w))
                begin
                    if(good[long_cpuid392/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid392 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid392/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid392])
        end // if (done[392])

        if (done[393]) begin
            timeout[long_cpuid393] = 0;
            //check_bad_trap(spc393_phy_pc_w, 393, long_cpuid393);
            if(active_thread[long_cpuid393])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc393_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid393/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 393 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid393]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc393_phy_pc_w))
                begin
                    if(good[long_cpuid393/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid393 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid393/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid393])
        end // if (done[393])

        if (done[394]) begin
            timeout[long_cpuid394] = 0;
            //check_bad_trap(spc394_phy_pc_w, 394, long_cpuid394);
            if(active_thread[long_cpuid394])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc394_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid394/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 394 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid394]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc394_phy_pc_w))
                begin
                    if(good[long_cpuid394/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid394 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid394/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid394])
        end // if (done[394])

        if (done[395]) begin
            timeout[long_cpuid395] = 0;
            //check_bad_trap(spc395_phy_pc_w, 395, long_cpuid395);
            if(active_thread[long_cpuid395])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc395_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid395/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 395 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid395]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc395_phy_pc_w))
                begin
                    if(good[long_cpuid395/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid395 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid395/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid395])
        end // if (done[395])

        if (done[396]) begin
            timeout[long_cpuid396] = 0;
            //check_bad_trap(spc396_phy_pc_w, 396, long_cpuid396);
            if(active_thread[long_cpuid396])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc396_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid396/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 396 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid396]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc396_phy_pc_w))
                begin
                    if(good[long_cpuid396/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid396 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid396/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid396])
        end // if (done[396])

        if (done[397]) begin
            timeout[long_cpuid397] = 0;
            //check_bad_trap(spc397_phy_pc_w, 397, long_cpuid397);
            if(active_thread[long_cpuid397])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc397_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid397/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 397 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid397]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc397_phy_pc_w))
                begin
                    if(good[long_cpuid397/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid397 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid397/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid397])
        end // if (done[397])

        if (done[398]) begin
            timeout[long_cpuid398] = 0;
            //check_bad_trap(spc398_phy_pc_w, 398, long_cpuid398);
            if(active_thread[long_cpuid398])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc398_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid398/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 398 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid398]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc398_phy_pc_w))
                begin
                    if(good[long_cpuid398/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid398 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid398/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid398])
        end // if (done[398])

        if (done[399]) begin
            timeout[long_cpuid399] = 0;
            //check_bad_trap(spc399_phy_pc_w, 399, long_cpuid399);
            if(active_thread[long_cpuid399])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc399_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid399/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 399 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid399]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc399_phy_pc_w))
                begin
                    if(good[long_cpuid399/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid399 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid399/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid399])
        end // if (done[399])

        if (done[400]) begin
            timeout[long_cpuid400] = 0;
            //check_bad_trap(spc400_phy_pc_w, 400, long_cpuid400);
            if(active_thread[long_cpuid400])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc400_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid400/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 400 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid400]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc400_phy_pc_w))
                begin
                    if(good[long_cpuid400/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid400 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid400/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid400])
        end // if (done[400])

        if (done[401]) begin
            timeout[long_cpuid401] = 0;
            //check_bad_trap(spc401_phy_pc_w, 401, long_cpuid401);
            if(active_thread[long_cpuid401])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc401_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid401/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 401 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid401]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc401_phy_pc_w))
                begin
                    if(good[long_cpuid401/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid401 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid401/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid401])
        end // if (done[401])

        if (done[402]) begin
            timeout[long_cpuid402] = 0;
            //check_bad_trap(spc402_phy_pc_w, 402, long_cpuid402);
            if(active_thread[long_cpuid402])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc402_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid402/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 402 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid402]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc402_phy_pc_w))
                begin
                    if(good[long_cpuid402/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid402 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid402/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid402])
        end // if (done[402])

        if (done[403]) begin
            timeout[long_cpuid403] = 0;
            //check_bad_trap(spc403_phy_pc_w, 403, long_cpuid403);
            if(active_thread[long_cpuid403])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc403_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid403/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 403 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid403]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc403_phy_pc_w))
                begin
                    if(good[long_cpuid403/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid403 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid403/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid403])
        end // if (done[403])

        if (done[404]) begin
            timeout[long_cpuid404] = 0;
            //check_bad_trap(spc404_phy_pc_w, 404, long_cpuid404);
            if(active_thread[long_cpuid404])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc404_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid404/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 404 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid404]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc404_phy_pc_w))
                begin
                    if(good[long_cpuid404/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid404 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid404/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid404])
        end // if (done[404])

        if (done[405]) begin
            timeout[long_cpuid405] = 0;
            //check_bad_trap(spc405_phy_pc_w, 405, long_cpuid405);
            if(active_thread[long_cpuid405])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc405_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid405/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 405 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid405]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc405_phy_pc_w))
                begin
                    if(good[long_cpuid405/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid405 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid405/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid405])
        end // if (done[405])

        if (done[406]) begin
            timeout[long_cpuid406] = 0;
            //check_bad_trap(spc406_phy_pc_w, 406, long_cpuid406);
            if(active_thread[long_cpuid406])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc406_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid406/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 406 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid406]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc406_phy_pc_w))
                begin
                    if(good[long_cpuid406/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid406 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid406/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid406])
        end // if (done[406])

        if (done[407]) begin
            timeout[long_cpuid407] = 0;
            //check_bad_trap(spc407_phy_pc_w, 407, long_cpuid407);
            if(active_thread[long_cpuid407])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc407_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid407/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 407 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid407]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc407_phy_pc_w))
                begin
                    if(good[long_cpuid407/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid407 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid407/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid407])
        end // if (done[407])

        if (done[408]) begin
            timeout[long_cpuid408] = 0;
            //check_bad_trap(spc408_phy_pc_w, 408, long_cpuid408);
            if(active_thread[long_cpuid408])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc408_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid408/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 408 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid408]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc408_phy_pc_w))
                begin
                    if(good[long_cpuid408/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid408 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid408/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid408])
        end // if (done[408])

        if (done[409]) begin
            timeout[long_cpuid409] = 0;
            //check_bad_trap(spc409_phy_pc_w, 409, long_cpuid409);
            if(active_thread[long_cpuid409])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc409_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid409/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 409 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid409]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc409_phy_pc_w))
                begin
                    if(good[long_cpuid409/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid409 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid409/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid409])
        end // if (done[409])

        if (done[410]) begin
            timeout[long_cpuid410] = 0;
            //check_bad_trap(spc410_phy_pc_w, 410, long_cpuid410);
            if(active_thread[long_cpuid410])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc410_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid410/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 410 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid410]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc410_phy_pc_w))
                begin
                    if(good[long_cpuid410/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid410 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid410/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid410])
        end // if (done[410])

        if (done[411]) begin
            timeout[long_cpuid411] = 0;
            //check_bad_trap(spc411_phy_pc_w, 411, long_cpuid411);
            if(active_thread[long_cpuid411])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc411_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid411/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 411 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid411]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc411_phy_pc_w))
                begin
                    if(good[long_cpuid411/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid411 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid411/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid411])
        end // if (done[411])

        if (done[412]) begin
            timeout[long_cpuid412] = 0;
            //check_bad_trap(spc412_phy_pc_w, 412, long_cpuid412);
            if(active_thread[long_cpuid412])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc412_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid412/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 412 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid412]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc412_phy_pc_w))
                begin
                    if(good[long_cpuid412/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid412 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid412/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid412])
        end // if (done[412])

        if (done[413]) begin
            timeout[long_cpuid413] = 0;
            //check_bad_trap(spc413_phy_pc_w, 413, long_cpuid413);
            if(active_thread[long_cpuid413])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc413_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid413/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 413 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid413]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc413_phy_pc_w))
                begin
                    if(good[long_cpuid413/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid413 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid413/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid413])
        end // if (done[413])

        if (done[414]) begin
            timeout[long_cpuid414] = 0;
            //check_bad_trap(spc414_phy_pc_w, 414, long_cpuid414);
            if(active_thread[long_cpuid414])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc414_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid414/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 414 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid414]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc414_phy_pc_w))
                begin
                    if(good[long_cpuid414/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid414 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid414/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid414])
        end // if (done[414])

        if (done[415]) begin
            timeout[long_cpuid415] = 0;
            //check_bad_trap(spc415_phy_pc_w, 415, long_cpuid415);
            if(active_thread[long_cpuid415])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc415_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid415/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 415 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid415]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc415_phy_pc_w))
                begin
                    if(good[long_cpuid415/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid415 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid415/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid415])
        end // if (done[415])

        if (done[416]) begin
            timeout[long_cpuid416] = 0;
            //check_bad_trap(spc416_phy_pc_w, 416, long_cpuid416);
            if(active_thread[long_cpuid416])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc416_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid416/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 416 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid416]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc416_phy_pc_w))
                begin
                    if(good[long_cpuid416/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid416 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid416/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid416])
        end // if (done[416])

        if (done[417]) begin
            timeout[long_cpuid417] = 0;
            //check_bad_trap(spc417_phy_pc_w, 417, long_cpuid417);
            if(active_thread[long_cpuid417])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc417_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid417/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 417 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid417]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc417_phy_pc_w))
                begin
                    if(good[long_cpuid417/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid417 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid417/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid417])
        end // if (done[417])

        if (done[418]) begin
            timeout[long_cpuid418] = 0;
            //check_bad_trap(spc418_phy_pc_w, 418, long_cpuid418);
            if(active_thread[long_cpuid418])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc418_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid418/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 418 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid418]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc418_phy_pc_w))
                begin
                    if(good[long_cpuid418/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid418 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid418/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid418])
        end // if (done[418])

        if (done[419]) begin
            timeout[long_cpuid419] = 0;
            //check_bad_trap(spc419_phy_pc_w, 419, long_cpuid419);
            if(active_thread[long_cpuid419])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc419_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid419/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 419 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid419]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc419_phy_pc_w))
                begin
                    if(good[long_cpuid419/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid419 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid419/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid419])
        end // if (done[419])

        if (done[420]) begin
            timeout[long_cpuid420] = 0;
            //check_bad_trap(spc420_phy_pc_w, 420, long_cpuid420);
            if(active_thread[long_cpuid420])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc420_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid420/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 420 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid420]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc420_phy_pc_w))
                begin
                    if(good[long_cpuid420/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid420 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid420/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid420])
        end // if (done[420])

        if (done[421]) begin
            timeout[long_cpuid421] = 0;
            //check_bad_trap(spc421_phy_pc_w, 421, long_cpuid421);
            if(active_thread[long_cpuid421])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc421_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid421/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 421 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid421]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc421_phy_pc_w))
                begin
                    if(good[long_cpuid421/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid421 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid421/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid421])
        end // if (done[421])

        if (done[422]) begin
            timeout[long_cpuid422] = 0;
            //check_bad_trap(spc422_phy_pc_w, 422, long_cpuid422);
            if(active_thread[long_cpuid422])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc422_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid422/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 422 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid422]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc422_phy_pc_w))
                begin
                    if(good[long_cpuid422/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid422 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid422/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid422])
        end // if (done[422])

        if (done[423]) begin
            timeout[long_cpuid423] = 0;
            //check_bad_trap(spc423_phy_pc_w, 423, long_cpuid423);
            if(active_thread[long_cpuid423])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc423_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid423/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 423 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid423]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc423_phy_pc_w))
                begin
                    if(good[long_cpuid423/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid423 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid423/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid423])
        end // if (done[423])

        if (done[424]) begin
            timeout[long_cpuid424] = 0;
            //check_bad_trap(spc424_phy_pc_w, 424, long_cpuid424);
            if(active_thread[long_cpuid424])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc424_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid424/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 424 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid424]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc424_phy_pc_w))
                begin
                    if(good[long_cpuid424/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid424 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid424/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid424])
        end // if (done[424])

        if (done[425]) begin
            timeout[long_cpuid425] = 0;
            //check_bad_trap(spc425_phy_pc_w, 425, long_cpuid425);
            if(active_thread[long_cpuid425])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc425_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid425/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 425 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid425]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc425_phy_pc_w))
                begin
                    if(good[long_cpuid425/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid425 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid425/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid425])
        end // if (done[425])

        if (done[426]) begin
            timeout[long_cpuid426] = 0;
            //check_bad_trap(spc426_phy_pc_w, 426, long_cpuid426);
            if(active_thread[long_cpuid426])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc426_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid426/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 426 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid426]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc426_phy_pc_w))
                begin
                    if(good[long_cpuid426/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid426 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid426/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid426])
        end // if (done[426])

        if (done[427]) begin
            timeout[long_cpuid427] = 0;
            //check_bad_trap(spc427_phy_pc_w, 427, long_cpuid427);
            if(active_thread[long_cpuid427])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc427_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid427/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 427 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid427]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc427_phy_pc_w))
                begin
                    if(good[long_cpuid427/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid427 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid427/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid427])
        end // if (done[427])

        if (done[428]) begin
            timeout[long_cpuid428] = 0;
            //check_bad_trap(spc428_phy_pc_w, 428, long_cpuid428);
            if(active_thread[long_cpuid428])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc428_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid428/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 428 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid428]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc428_phy_pc_w))
                begin
                    if(good[long_cpuid428/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid428 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid428/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid428])
        end // if (done[428])

        if (done[429]) begin
            timeout[long_cpuid429] = 0;
            //check_bad_trap(spc429_phy_pc_w, 429, long_cpuid429);
            if(active_thread[long_cpuid429])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc429_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid429/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 429 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid429]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc429_phy_pc_w))
                begin
                    if(good[long_cpuid429/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid429 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid429/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid429])
        end // if (done[429])

        if (done[430]) begin
            timeout[long_cpuid430] = 0;
            //check_bad_trap(spc430_phy_pc_w, 430, long_cpuid430);
            if(active_thread[long_cpuid430])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc430_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid430/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 430 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid430]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc430_phy_pc_w))
                begin
                    if(good[long_cpuid430/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid430 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid430/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid430])
        end // if (done[430])

        if (done[431]) begin
            timeout[long_cpuid431] = 0;
            //check_bad_trap(spc431_phy_pc_w, 431, long_cpuid431);
            if(active_thread[long_cpuid431])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc431_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid431/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 431 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid431]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc431_phy_pc_w))
                begin
                    if(good[long_cpuid431/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid431 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid431/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid431])
        end // if (done[431])

        if (done[432]) begin
            timeout[long_cpuid432] = 0;
            //check_bad_trap(spc432_phy_pc_w, 432, long_cpuid432);
            if(active_thread[long_cpuid432])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc432_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid432/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 432 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid432]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc432_phy_pc_w))
                begin
                    if(good[long_cpuid432/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid432 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid432/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid432])
        end // if (done[432])

        if (done[433]) begin
            timeout[long_cpuid433] = 0;
            //check_bad_trap(spc433_phy_pc_w, 433, long_cpuid433);
            if(active_thread[long_cpuid433])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc433_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid433/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 433 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid433]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc433_phy_pc_w))
                begin
                    if(good[long_cpuid433/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid433 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid433/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid433])
        end // if (done[433])

        if (done[434]) begin
            timeout[long_cpuid434] = 0;
            //check_bad_trap(spc434_phy_pc_w, 434, long_cpuid434);
            if(active_thread[long_cpuid434])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc434_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid434/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 434 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid434]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc434_phy_pc_w))
                begin
                    if(good[long_cpuid434/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid434 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid434/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid434])
        end // if (done[434])

        if (done[435]) begin
            timeout[long_cpuid435] = 0;
            //check_bad_trap(spc435_phy_pc_w, 435, long_cpuid435);
            if(active_thread[long_cpuid435])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc435_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid435/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 435 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid435]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc435_phy_pc_w))
                begin
                    if(good[long_cpuid435/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid435 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid435/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid435])
        end // if (done[435])

        if (done[436]) begin
            timeout[long_cpuid436] = 0;
            //check_bad_trap(spc436_phy_pc_w, 436, long_cpuid436);
            if(active_thread[long_cpuid436])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc436_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid436/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 436 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid436]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc436_phy_pc_w))
                begin
                    if(good[long_cpuid436/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid436 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid436/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid436])
        end // if (done[436])

        if (done[437]) begin
            timeout[long_cpuid437] = 0;
            //check_bad_trap(spc437_phy_pc_w, 437, long_cpuid437);
            if(active_thread[long_cpuid437])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc437_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid437/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 437 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid437]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc437_phy_pc_w))
                begin
                    if(good[long_cpuid437/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid437 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid437/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid437])
        end // if (done[437])

        if (done[438]) begin
            timeout[long_cpuid438] = 0;
            //check_bad_trap(spc438_phy_pc_w, 438, long_cpuid438);
            if(active_thread[long_cpuid438])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc438_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid438/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 438 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid438]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc438_phy_pc_w))
                begin
                    if(good[long_cpuid438/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid438 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid438/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid438])
        end // if (done[438])

        if (done[439]) begin
            timeout[long_cpuid439] = 0;
            //check_bad_trap(spc439_phy_pc_w, 439, long_cpuid439);
            if(active_thread[long_cpuid439])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc439_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid439/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 439 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid439]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc439_phy_pc_w))
                begin
                    if(good[long_cpuid439/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid439 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid439/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid439])
        end // if (done[439])

        if (done[440]) begin
            timeout[long_cpuid440] = 0;
            //check_bad_trap(spc440_phy_pc_w, 440, long_cpuid440);
            if(active_thread[long_cpuid440])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc440_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid440/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 440 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid440]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc440_phy_pc_w))
                begin
                    if(good[long_cpuid440/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid440 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid440/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid440])
        end // if (done[440])

        if (done[441]) begin
            timeout[long_cpuid441] = 0;
            //check_bad_trap(spc441_phy_pc_w, 441, long_cpuid441);
            if(active_thread[long_cpuid441])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc441_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid441/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 441 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid441]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc441_phy_pc_w))
                begin
                    if(good[long_cpuid441/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid441 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid441/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid441])
        end // if (done[441])

        if (done[442]) begin
            timeout[long_cpuid442] = 0;
            //check_bad_trap(spc442_phy_pc_w, 442, long_cpuid442);
            if(active_thread[long_cpuid442])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc442_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid442/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 442 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid442]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc442_phy_pc_w))
                begin
                    if(good[long_cpuid442/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid442 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid442/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid442])
        end // if (done[442])

        if (done[443]) begin
            timeout[long_cpuid443] = 0;
            //check_bad_trap(spc443_phy_pc_w, 443, long_cpuid443);
            if(active_thread[long_cpuid443])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc443_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid443/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 443 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid443]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc443_phy_pc_w))
                begin
                    if(good[long_cpuid443/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid443 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid443/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid443])
        end // if (done[443])

        if (done[444]) begin
            timeout[long_cpuid444] = 0;
            //check_bad_trap(spc444_phy_pc_w, 444, long_cpuid444);
            if(active_thread[long_cpuid444])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc444_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid444/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 444 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid444]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc444_phy_pc_w))
                begin
                    if(good[long_cpuid444/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid444 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid444/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid444])
        end // if (done[444])

        if (done[445]) begin
            timeout[long_cpuid445] = 0;
            //check_bad_trap(spc445_phy_pc_w, 445, long_cpuid445);
            if(active_thread[long_cpuid445])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc445_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid445/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 445 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid445]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc445_phy_pc_w))
                begin
                    if(good[long_cpuid445/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid445 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid445/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid445])
        end // if (done[445])

        if (done[446]) begin
            timeout[long_cpuid446] = 0;
            //check_bad_trap(spc446_phy_pc_w, 446, long_cpuid446);
            if(active_thread[long_cpuid446])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc446_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid446/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 446 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid446]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc446_phy_pc_w))
                begin
                    if(good[long_cpuid446/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid446 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid446/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid446])
        end // if (done[446])

        if (done[447]) begin
            timeout[long_cpuid447] = 0;
            //check_bad_trap(spc447_phy_pc_w, 447, long_cpuid447);
            if(active_thread[long_cpuid447])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc447_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid447/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 447 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid447]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc447_phy_pc_w))
                begin
                    if(good[long_cpuid447/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid447 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid447/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid447])
        end // if (done[447])

        if (done[448]) begin
            timeout[long_cpuid448] = 0;
            //check_bad_trap(spc448_phy_pc_w, 448, long_cpuid448);
            if(active_thread[long_cpuid448])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc448_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid448/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 448 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid448]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc448_phy_pc_w))
                begin
                    if(good[long_cpuid448/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid448 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid448/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid448])
        end // if (done[448])

        if (done[449]) begin
            timeout[long_cpuid449] = 0;
            //check_bad_trap(spc449_phy_pc_w, 449, long_cpuid449);
            if(active_thread[long_cpuid449])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc449_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid449/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 449 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid449]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc449_phy_pc_w))
                begin
                    if(good[long_cpuid449/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid449 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid449/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid449])
        end // if (done[449])

        if (done[450]) begin
            timeout[long_cpuid450] = 0;
            //check_bad_trap(spc450_phy_pc_w, 450, long_cpuid450);
            if(active_thread[long_cpuid450])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc450_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid450/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 450 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid450]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc450_phy_pc_w))
                begin
                    if(good[long_cpuid450/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid450 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid450/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid450])
        end // if (done[450])

        if (done[451]) begin
            timeout[long_cpuid451] = 0;
            //check_bad_trap(spc451_phy_pc_w, 451, long_cpuid451);
            if(active_thread[long_cpuid451])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc451_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid451/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 451 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid451]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc451_phy_pc_w))
                begin
                    if(good[long_cpuid451/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid451 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid451/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid451])
        end // if (done[451])

        if (done[452]) begin
            timeout[long_cpuid452] = 0;
            //check_bad_trap(spc452_phy_pc_w, 452, long_cpuid452);
            if(active_thread[long_cpuid452])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc452_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid452/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 452 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid452]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc452_phy_pc_w))
                begin
                    if(good[long_cpuid452/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid452 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid452/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid452])
        end // if (done[452])

        if (done[453]) begin
            timeout[long_cpuid453] = 0;
            //check_bad_trap(spc453_phy_pc_w, 453, long_cpuid453);
            if(active_thread[long_cpuid453])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc453_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid453/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 453 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid453]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc453_phy_pc_w))
                begin
                    if(good[long_cpuid453/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid453 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid453/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid453])
        end // if (done[453])

        if (done[454]) begin
            timeout[long_cpuid454] = 0;
            //check_bad_trap(spc454_phy_pc_w, 454, long_cpuid454);
            if(active_thread[long_cpuid454])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc454_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid454/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 454 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid454]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc454_phy_pc_w))
                begin
                    if(good[long_cpuid454/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid454 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid454/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid454])
        end // if (done[454])

        if (done[455]) begin
            timeout[long_cpuid455] = 0;
            //check_bad_trap(spc455_phy_pc_w, 455, long_cpuid455);
            if(active_thread[long_cpuid455])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc455_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid455/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 455 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid455]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc455_phy_pc_w))
                begin
                    if(good[long_cpuid455/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid455 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid455/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid455])
        end // if (done[455])

        if (done[456]) begin
            timeout[long_cpuid456] = 0;
            //check_bad_trap(spc456_phy_pc_w, 456, long_cpuid456);
            if(active_thread[long_cpuid456])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc456_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid456/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 456 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid456]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc456_phy_pc_w))
                begin
                    if(good[long_cpuid456/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid456 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid456/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid456])
        end // if (done[456])

        if (done[457]) begin
            timeout[long_cpuid457] = 0;
            //check_bad_trap(spc457_phy_pc_w, 457, long_cpuid457);
            if(active_thread[long_cpuid457])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc457_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid457/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 457 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid457]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc457_phy_pc_w))
                begin
                    if(good[long_cpuid457/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid457 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid457/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid457])
        end // if (done[457])

        if (done[458]) begin
            timeout[long_cpuid458] = 0;
            //check_bad_trap(spc458_phy_pc_w, 458, long_cpuid458);
            if(active_thread[long_cpuid458])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc458_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid458/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 458 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid458]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc458_phy_pc_w))
                begin
                    if(good[long_cpuid458/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid458 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid458/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid458])
        end // if (done[458])

        if (done[459]) begin
            timeout[long_cpuid459] = 0;
            //check_bad_trap(spc459_phy_pc_w, 459, long_cpuid459);
            if(active_thread[long_cpuid459])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc459_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid459/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 459 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid459]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc459_phy_pc_w))
                begin
                    if(good[long_cpuid459/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid459 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid459/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid459])
        end // if (done[459])

        if (done[460]) begin
            timeout[long_cpuid460] = 0;
            //check_bad_trap(spc460_phy_pc_w, 460, long_cpuid460);
            if(active_thread[long_cpuid460])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc460_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid460/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 460 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid460]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc460_phy_pc_w))
                begin
                    if(good[long_cpuid460/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid460 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid460/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid460])
        end // if (done[460])

        if (done[461]) begin
            timeout[long_cpuid461] = 0;
            //check_bad_trap(spc461_phy_pc_w, 461, long_cpuid461);
            if(active_thread[long_cpuid461])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc461_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid461/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 461 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid461]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc461_phy_pc_w))
                begin
                    if(good[long_cpuid461/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid461 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid461/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid461])
        end // if (done[461])

        if (done[462]) begin
            timeout[long_cpuid462] = 0;
            //check_bad_trap(spc462_phy_pc_w, 462, long_cpuid462);
            if(active_thread[long_cpuid462])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc462_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid462/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 462 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid462]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc462_phy_pc_w))
                begin
                    if(good[long_cpuid462/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid462 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid462/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid462])
        end // if (done[462])

        if (done[463]) begin
            timeout[long_cpuid463] = 0;
            //check_bad_trap(spc463_phy_pc_w, 463, long_cpuid463);
            if(active_thread[long_cpuid463])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc463_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid463/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 463 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid463]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc463_phy_pc_w))
                begin
                    if(good[long_cpuid463/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid463 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid463/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid463])
        end // if (done[463])

        if (done[464]) begin
            timeout[long_cpuid464] = 0;
            //check_bad_trap(spc464_phy_pc_w, 464, long_cpuid464);
            if(active_thread[long_cpuid464])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc464_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid464/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 464 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid464]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc464_phy_pc_w))
                begin
                    if(good[long_cpuid464/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid464 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid464/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid464])
        end // if (done[464])

        if (done[465]) begin
            timeout[long_cpuid465] = 0;
            //check_bad_trap(spc465_phy_pc_w, 465, long_cpuid465);
            if(active_thread[long_cpuid465])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc465_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid465/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 465 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid465]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc465_phy_pc_w))
                begin
                    if(good[long_cpuid465/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid465 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid465/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid465])
        end // if (done[465])

        if (done[466]) begin
            timeout[long_cpuid466] = 0;
            //check_bad_trap(spc466_phy_pc_w, 466, long_cpuid466);
            if(active_thread[long_cpuid466])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc466_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid466/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 466 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid466]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc466_phy_pc_w))
                begin
                    if(good[long_cpuid466/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid466 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid466/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid466])
        end // if (done[466])

        if (done[467]) begin
            timeout[long_cpuid467] = 0;
            //check_bad_trap(spc467_phy_pc_w, 467, long_cpuid467);
            if(active_thread[long_cpuid467])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc467_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid467/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 467 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid467]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc467_phy_pc_w))
                begin
                    if(good[long_cpuid467/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid467 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid467/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid467])
        end // if (done[467])

        if (done[468]) begin
            timeout[long_cpuid468] = 0;
            //check_bad_trap(spc468_phy_pc_w, 468, long_cpuid468);
            if(active_thread[long_cpuid468])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc468_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid468/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 468 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid468]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc468_phy_pc_w))
                begin
                    if(good[long_cpuid468/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid468 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid468/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid468])
        end // if (done[468])

        if (done[469]) begin
            timeout[long_cpuid469] = 0;
            //check_bad_trap(spc469_phy_pc_w, 469, long_cpuid469);
            if(active_thread[long_cpuid469])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc469_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid469/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 469 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid469]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc469_phy_pc_w))
                begin
                    if(good[long_cpuid469/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid469 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid469/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid469])
        end // if (done[469])

        if (done[470]) begin
            timeout[long_cpuid470] = 0;
            //check_bad_trap(spc470_phy_pc_w, 470, long_cpuid470);
            if(active_thread[long_cpuid470])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc470_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid470/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 470 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid470]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc470_phy_pc_w))
                begin
                    if(good[long_cpuid470/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid470 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid470/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid470])
        end // if (done[470])

        if (done[471]) begin
            timeout[long_cpuid471] = 0;
            //check_bad_trap(spc471_phy_pc_w, 471, long_cpuid471);
            if(active_thread[long_cpuid471])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc471_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid471/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 471 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid471]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc471_phy_pc_w))
                begin
                    if(good[long_cpuid471/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid471 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid471/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid471])
        end // if (done[471])

        if (done[472]) begin
            timeout[long_cpuid472] = 0;
            //check_bad_trap(spc472_phy_pc_w, 472, long_cpuid472);
            if(active_thread[long_cpuid472])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc472_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid472/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 472 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid472]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc472_phy_pc_w))
                begin
                    if(good[long_cpuid472/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid472 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid472/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid472])
        end // if (done[472])

        if (done[473]) begin
            timeout[long_cpuid473] = 0;
            //check_bad_trap(spc473_phy_pc_w, 473, long_cpuid473);
            if(active_thread[long_cpuid473])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc473_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid473/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 473 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid473]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc473_phy_pc_w))
                begin
                    if(good[long_cpuid473/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid473 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid473/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid473])
        end // if (done[473])

        if (done[474]) begin
            timeout[long_cpuid474] = 0;
            //check_bad_trap(spc474_phy_pc_w, 474, long_cpuid474);
            if(active_thread[long_cpuid474])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc474_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid474/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 474 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid474]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc474_phy_pc_w))
                begin
                    if(good[long_cpuid474/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid474 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid474/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid474])
        end // if (done[474])

        if (done[475]) begin
            timeout[long_cpuid475] = 0;
            //check_bad_trap(spc475_phy_pc_w, 475, long_cpuid475);
            if(active_thread[long_cpuid475])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc475_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid475/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 475 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid475]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc475_phy_pc_w))
                begin
                    if(good[long_cpuid475/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid475 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid475/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid475])
        end // if (done[475])

        if (done[476]) begin
            timeout[long_cpuid476] = 0;
            //check_bad_trap(spc476_phy_pc_w, 476, long_cpuid476);
            if(active_thread[long_cpuid476])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc476_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid476/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 476 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid476]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc476_phy_pc_w))
                begin
                    if(good[long_cpuid476/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid476 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid476/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid476])
        end // if (done[476])

        if (done[477]) begin
            timeout[long_cpuid477] = 0;
            //check_bad_trap(spc477_phy_pc_w, 477, long_cpuid477);
            if(active_thread[long_cpuid477])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc477_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid477/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 477 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid477]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc477_phy_pc_w))
                begin
                    if(good[long_cpuid477/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid477 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid477/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid477])
        end // if (done[477])

        if (done[478]) begin
            timeout[long_cpuid478] = 0;
            //check_bad_trap(spc478_phy_pc_w, 478, long_cpuid478);
            if(active_thread[long_cpuid478])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc478_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid478/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 478 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid478]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc478_phy_pc_w))
                begin
                    if(good[long_cpuid478/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid478 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid478/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid478])
        end // if (done[478])

        if (done[479]) begin
            timeout[long_cpuid479] = 0;
            //check_bad_trap(spc479_phy_pc_w, 479, long_cpuid479);
            if(active_thread[long_cpuid479])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc479_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid479/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 479 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid479]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc479_phy_pc_w))
                begin
                    if(good[long_cpuid479/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid479 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid479/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid479])
        end // if (done[479])

        if (done[480]) begin
            timeout[long_cpuid480] = 0;
            //check_bad_trap(spc480_phy_pc_w, 480, long_cpuid480);
            if(active_thread[long_cpuid480])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc480_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid480/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 480 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid480]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc480_phy_pc_w))
                begin
                    if(good[long_cpuid480/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid480 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid480/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid480])
        end // if (done[480])

        if (done[481]) begin
            timeout[long_cpuid481] = 0;
            //check_bad_trap(spc481_phy_pc_w, 481, long_cpuid481);
            if(active_thread[long_cpuid481])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc481_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid481/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 481 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid481]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc481_phy_pc_w))
                begin
                    if(good[long_cpuid481/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid481 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid481/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid481])
        end // if (done[481])

        if (done[482]) begin
            timeout[long_cpuid482] = 0;
            //check_bad_trap(spc482_phy_pc_w, 482, long_cpuid482);
            if(active_thread[long_cpuid482])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc482_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid482/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 482 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid482]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc482_phy_pc_w))
                begin
                    if(good[long_cpuid482/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid482 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid482/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid482])
        end // if (done[482])

        if (done[483]) begin
            timeout[long_cpuid483] = 0;
            //check_bad_trap(spc483_phy_pc_w, 483, long_cpuid483);
            if(active_thread[long_cpuid483])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc483_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid483/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 483 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid483]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc483_phy_pc_w))
                begin
                    if(good[long_cpuid483/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid483 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid483/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid483])
        end // if (done[483])

        if (done[484]) begin
            timeout[long_cpuid484] = 0;
            //check_bad_trap(spc484_phy_pc_w, 484, long_cpuid484);
            if(active_thread[long_cpuid484])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc484_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid484/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 484 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid484]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc484_phy_pc_w))
                begin
                    if(good[long_cpuid484/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid484 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid484/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid484])
        end // if (done[484])

        if (done[485]) begin
            timeout[long_cpuid485] = 0;
            //check_bad_trap(spc485_phy_pc_w, 485, long_cpuid485);
            if(active_thread[long_cpuid485])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc485_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid485/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 485 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid485]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc485_phy_pc_w))
                begin
                    if(good[long_cpuid485/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid485 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid485/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid485])
        end // if (done[485])

        if (done[486]) begin
            timeout[long_cpuid486] = 0;
            //check_bad_trap(spc486_phy_pc_w, 486, long_cpuid486);
            if(active_thread[long_cpuid486])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc486_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid486/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 486 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid486]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc486_phy_pc_w))
                begin
                    if(good[long_cpuid486/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid486 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid486/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid486])
        end // if (done[486])

        if (done[487]) begin
            timeout[long_cpuid487] = 0;
            //check_bad_trap(spc487_phy_pc_w, 487, long_cpuid487);
            if(active_thread[long_cpuid487])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc487_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid487/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 487 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid487]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc487_phy_pc_w))
                begin
                    if(good[long_cpuid487/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid487 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid487/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid487])
        end // if (done[487])

        if (done[488]) begin
            timeout[long_cpuid488] = 0;
            //check_bad_trap(spc488_phy_pc_w, 488, long_cpuid488);
            if(active_thread[long_cpuid488])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc488_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid488/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 488 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid488]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc488_phy_pc_w))
                begin
                    if(good[long_cpuid488/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid488 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid488/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid488])
        end // if (done[488])

        if (done[489]) begin
            timeout[long_cpuid489] = 0;
            //check_bad_trap(spc489_phy_pc_w, 489, long_cpuid489);
            if(active_thread[long_cpuid489])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc489_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid489/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 489 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid489]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc489_phy_pc_w))
                begin
                    if(good[long_cpuid489/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid489 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid489/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid489])
        end // if (done[489])

        if (done[490]) begin
            timeout[long_cpuid490] = 0;
            //check_bad_trap(spc490_phy_pc_w, 490, long_cpuid490);
            if(active_thread[long_cpuid490])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc490_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid490/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 490 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid490]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc490_phy_pc_w))
                begin
                    if(good[long_cpuid490/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid490 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid490/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid490])
        end // if (done[490])

        if (done[491]) begin
            timeout[long_cpuid491] = 0;
            //check_bad_trap(spc491_phy_pc_w, 491, long_cpuid491);
            if(active_thread[long_cpuid491])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc491_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid491/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 491 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid491]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc491_phy_pc_w))
                begin
                    if(good[long_cpuid491/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid491 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid491/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid491])
        end // if (done[491])

        if (done[492]) begin
            timeout[long_cpuid492] = 0;
            //check_bad_trap(spc492_phy_pc_w, 492, long_cpuid492);
            if(active_thread[long_cpuid492])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc492_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid492/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 492 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid492]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc492_phy_pc_w))
                begin
                    if(good[long_cpuid492/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid492 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid492/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid492])
        end // if (done[492])

        if (done[493]) begin
            timeout[long_cpuid493] = 0;
            //check_bad_trap(spc493_phy_pc_w, 493, long_cpuid493);
            if(active_thread[long_cpuid493])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc493_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid493/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 493 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid493]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc493_phy_pc_w))
                begin
                    if(good[long_cpuid493/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid493 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid493/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid493])
        end // if (done[493])

        if (done[494]) begin
            timeout[long_cpuid494] = 0;
            //check_bad_trap(spc494_phy_pc_w, 494, long_cpuid494);
            if(active_thread[long_cpuid494])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc494_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid494/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 494 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid494]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc494_phy_pc_w))
                begin
                    if(good[long_cpuid494/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid494 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid494/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid494])
        end // if (done[494])

        if (done[495]) begin
            timeout[long_cpuid495] = 0;
            //check_bad_trap(spc495_phy_pc_w, 495, long_cpuid495);
            if(active_thread[long_cpuid495])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc495_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid495/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 495 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid495]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc495_phy_pc_w))
                begin
                    if(good[long_cpuid495/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid495 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid495/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid495])
        end // if (done[495])

        if (done[496]) begin
            timeout[long_cpuid496] = 0;
            //check_bad_trap(spc496_phy_pc_w, 496, long_cpuid496);
            if(active_thread[long_cpuid496])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc496_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid496/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 496 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid496]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc496_phy_pc_w))
                begin
                    if(good[long_cpuid496/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid496 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid496/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid496])
        end // if (done[496])

        if (done[497]) begin
            timeout[long_cpuid497] = 0;
            //check_bad_trap(spc497_phy_pc_w, 497, long_cpuid497);
            if(active_thread[long_cpuid497])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc497_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid497/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 497 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid497]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc497_phy_pc_w))
                begin
                    if(good[long_cpuid497/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid497 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid497/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid497])
        end // if (done[497])

        if (done[498]) begin
            timeout[long_cpuid498] = 0;
            //check_bad_trap(spc498_phy_pc_w, 498, long_cpuid498);
            if(active_thread[long_cpuid498])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc498_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid498/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 498 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid498]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc498_phy_pc_w))
                begin
                    if(good[long_cpuid498/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid498 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid498/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid498])
        end // if (done[498])

        if (done[499]) begin
            timeout[long_cpuid499] = 0;
            //check_bad_trap(spc499_phy_pc_w, 499, long_cpuid499);
            if(active_thread[long_cpuid499])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc499_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid499/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 499 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid499]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc499_phy_pc_w))
                begin
                    if(good[long_cpuid499/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid499 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid499/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid499])
        end // if (done[499])

        if (done[500]) begin
            timeout[long_cpuid500] = 0;
            //check_bad_trap(spc500_phy_pc_w, 500, long_cpuid500);
            if(active_thread[long_cpuid500])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc500_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid500/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 500 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid500]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc500_phy_pc_w))
                begin
                    if(good[long_cpuid500/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid500 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid500/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid500])
        end // if (done[500])

        if (done[501]) begin
            timeout[long_cpuid501] = 0;
            //check_bad_trap(spc501_phy_pc_w, 501, long_cpuid501);
            if(active_thread[long_cpuid501])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc501_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid501/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 501 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid501]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc501_phy_pc_w))
                begin
                    if(good[long_cpuid501/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid501 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid501/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid501])
        end // if (done[501])

        if (done[502]) begin
            timeout[long_cpuid502] = 0;
            //check_bad_trap(spc502_phy_pc_w, 502, long_cpuid502);
            if(active_thread[long_cpuid502])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc502_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid502/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 502 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid502]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc502_phy_pc_w))
                begin
                    if(good[long_cpuid502/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid502 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid502/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid502])
        end // if (done[502])

        if (done[503]) begin
            timeout[long_cpuid503] = 0;
            //check_bad_trap(spc503_phy_pc_w, 503, long_cpuid503);
            if(active_thread[long_cpuid503])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc503_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid503/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 503 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid503]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc503_phy_pc_w))
                begin
                    if(good[long_cpuid503/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid503 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid503/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid503])
        end // if (done[503])

        if (done[504]) begin
            timeout[long_cpuid504] = 0;
            //check_bad_trap(spc504_phy_pc_w, 504, long_cpuid504);
            if(active_thread[long_cpuid504])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc504_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid504/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 504 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid504]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc504_phy_pc_w))
                begin
                    if(good[long_cpuid504/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid504 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid504/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid504])
        end // if (done[504])

        if (done[505]) begin
            timeout[long_cpuid505] = 0;
            //check_bad_trap(spc505_phy_pc_w, 505, long_cpuid505);
            if(active_thread[long_cpuid505])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc505_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid505/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 505 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid505]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc505_phy_pc_w))
                begin
                    if(good[long_cpuid505/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid505 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid505/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid505])
        end // if (done[505])

        if (done[506]) begin
            timeout[long_cpuid506] = 0;
            //check_bad_trap(spc506_phy_pc_w, 506, long_cpuid506);
            if(active_thread[long_cpuid506])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc506_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid506/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 506 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid506]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc506_phy_pc_w))
                begin
                    if(good[long_cpuid506/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid506 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid506/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid506])
        end // if (done[506])

        if (done[507]) begin
            timeout[long_cpuid507] = 0;
            //check_bad_trap(spc507_phy_pc_w, 507, long_cpuid507);
            if(active_thread[long_cpuid507])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc507_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid507/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 507 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid507]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc507_phy_pc_w))
                begin
                    if(good[long_cpuid507/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid507 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid507/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid507])
        end // if (done[507])

        if (done[508]) begin
            timeout[long_cpuid508] = 0;
            //check_bad_trap(spc508_phy_pc_w, 508, long_cpuid508);
            if(active_thread[long_cpuid508])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc508_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid508/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 508 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid508]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc508_phy_pc_w))
                begin
                    if(good[long_cpuid508/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid508 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid508/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid508])
        end // if (done[508])

        if (done[509]) begin
            timeout[long_cpuid509] = 0;
            //check_bad_trap(spc509_phy_pc_w, 509, long_cpuid509);
            if(active_thread[long_cpuid509])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc509_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid509/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 509 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid509]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc509_phy_pc_w))
                begin
                    if(good[long_cpuid509/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid509 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid509/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid509])
        end // if (done[509])

        if (done[510]) begin
            timeout[long_cpuid510] = 0;
            //check_bad_trap(spc510_phy_pc_w, 510, long_cpuid510);
            if(active_thread[long_cpuid510])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc510_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid510/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 510 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid510]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc510_phy_pc_w))
                begin
                    if(good[long_cpuid510/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid510 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid510/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid510])
        end // if (done[510])

        if (done[511]) begin
            timeout[long_cpuid511] = 0;
            //check_bad_trap(spc511_phy_pc_w, 511, long_cpuid511);
            if(active_thread[long_cpuid511])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc511_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid511/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 511 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid511]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc511_phy_pc_w))
                begin
                    if(good[long_cpuid511/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid511 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid511/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid511])
        end // if (done[511])

        if (done[512]) begin
            timeout[long_cpuid512] = 0;
            //check_bad_trap(spc512_phy_pc_w, 512, long_cpuid512);
            if(active_thread[long_cpuid512])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc512_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid512/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 512 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid512]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc512_phy_pc_w))
                begin
                    if(good[long_cpuid512/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid512 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid512/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid512])
        end // if (done[512])

        if (done[513]) begin
            timeout[long_cpuid513] = 0;
            //check_bad_trap(spc513_phy_pc_w, 513, long_cpuid513);
            if(active_thread[long_cpuid513])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc513_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid513/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 513 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid513]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc513_phy_pc_w))
                begin
                    if(good[long_cpuid513/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid513 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid513/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid513])
        end // if (done[513])

        if (done[514]) begin
            timeout[long_cpuid514] = 0;
            //check_bad_trap(spc514_phy_pc_w, 514, long_cpuid514);
            if(active_thread[long_cpuid514])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc514_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid514/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 514 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid514]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc514_phy_pc_w))
                begin
                    if(good[long_cpuid514/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid514 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid514/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid514])
        end // if (done[514])

        if (done[515]) begin
            timeout[long_cpuid515] = 0;
            //check_bad_trap(spc515_phy_pc_w, 515, long_cpuid515);
            if(active_thread[long_cpuid515])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc515_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid515/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 515 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid515]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc515_phy_pc_w))
                begin
                    if(good[long_cpuid515/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid515 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid515/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid515])
        end // if (done[515])

        if (done[516]) begin
            timeout[long_cpuid516] = 0;
            //check_bad_trap(spc516_phy_pc_w, 516, long_cpuid516);
            if(active_thread[long_cpuid516])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc516_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid516/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 516 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid516]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc516_phy_pc_w))
                begin
                    if(good[long_cpuid516/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid516 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid516/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid516])
        end // if (done[516])

        if (done[517]) begin
            timeout[long_cpuid517] = 0;
            //check_bad_trap(spc517_phy_pc_w, 517, long_cpuid517);
            if(active_thread[long_cpuid517])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc517_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid517/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 517 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid517]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc517_phy_pc_w))
                begin
                    if(good[long_cpuid517/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid517 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid517/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid517])
        end // if (done[517])

        if (done[518]) begin
            timeout[long_cpuid518] = 0;
            //check_bad_trap(spc518_phy_pc_w, 518, long_cpuid518);
            if(active_thread[long_cpuid518])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc518_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid518/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 518 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid518]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc518_phy_pc_w))
                begin
                    if(good[long_cpuid518/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid518 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid518/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid518])
        end // if (done[518])

        if (done[519]) begin
            timeout[long_cpuid519] = 0;
            //check_bad_trap(spc519_phy_pc_w, 519, long_cpuid519);
            if(active_thread[long_cpuid519])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc519_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid519/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 519 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid519]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc519_phy_pc_w))
                begin
                    if(good[long_cpuid519/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid519 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid519/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid519])
        end // if (done[519])

        if (done[520]) begin
            timeout[long_cpuid520] = 0;
            //check_bad_trap(spc520_phy_pc_w, 520, long_cpuid520);
            if(active_thread[long_cpuid520])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc520_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid520/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 520 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid520]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc520_phy_pc_w))
                begin
                    if(good[long_cpuid520/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid520 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid520/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid520])
        end // if (done[520])

        if (done[521]) begin
            timeout[long_cpuid521] = 0;
            //check_bad_trap(spc521_phy_pc_w, 521, long_cpuid521);
            if(active_thread[long_cpuid521])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc521_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid521/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 521 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid521]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc521_phy_pc_w))
                begin
                    if(good[long_cpuid521/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid521 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid521/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid521])
        end // if (done[521])

        if (done[522]) begin
            timeout[long_cpuid522] = 0;
            //check_bad_trap(spc522_phy_pc_w, 522, long_cpuid522);
            if(active_thread[long_cpuid522])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc522_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid522/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 522 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid522]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc522_phy_pc_w))
                begin
                    if(good[long_cpuid522/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid522 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid522/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid522])
        end // if (done[522])

        if (done[523]) begin
            timeout[long_cpuid523] = 0;
            //check_bad_trap(spc523_phy_pc_w, 523, long_cpuid523);
            if(active_thread[long_cpuid523])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc523_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid523/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 523 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid523]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc523_phy_pc_w))
                begin
                    if(good[long_cpuid523/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid523 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid523/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid523])
        end // if (done[523])

        if (done[524]) begin
            timeout[long_cpuid524] = 0;
            //check_bad_trap(spc524_phy_pc_w, 524, long_cpuid524);
            if(active_thread[long_cpuid524])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc524_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid524/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 524 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid524]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc524_phy_pc_w))
                begin
                    if(good[long_cpuid524/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid524 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid524/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid524])
        end // if (done[524])

        if (done[525]) begin
            timeout[long_cpuid525] = 0;
            //check_bad_trap(spc525_phy_pc_w, 525, long_cpuid525);
            if(active_thread[long_cpuid525])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc525_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid525/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 525 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid525]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc525_phy_pc_w))
                begin
                    if(good[long_cpuid525/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid525 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid525/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid525])
        end // if (done[525])

        if (done[526]) begin
            timeout[long_cpuid526] = 0;
            //check_bad_trap(spc526_phy_pc_w, 526, long_cpuid526);
            if(active_thread[long_cpuid526])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc526_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid526/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 526 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid526]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc526_phy_pc_w))
                begin
                    if(good[long_cpuid526/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid526 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid526/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid526])
        end // if (done[526])

        if (done[527]) begin
            timeout[long_cpuid527] = 0;
            //check_bad_trap(spc527_phy_pc_w, 527, long_cpuid527);
            if(active_thread[long_cpuid527])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc527_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid527/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 527 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid527]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc527_phy_pc_w))
                begin
                    if(good[long_cpuid527/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid527 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid527/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid527])
        end // if (done[527])

        if (done[528]) begin
            timeout[long_cpuid528] = 0;
            //check_bad_trap(spc528_phy_pc_w, 528, long_cpuid528);
            if(active_thread[long_cpuid528])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc528_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid528/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 528 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid528]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc528_phy_pc_w))
                begin
                    if(good[long_cpuid528/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid528 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid528/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid528])
        end // if (done[528])

        if (done[529]) begin
            timeout[long_cpuid529] = 0;
            //check_bad_trap(spc529_phy_pc_w, 529, long_cpuid529);
            if(active_thread[long_cpuid529])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc529_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid529/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 529 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid529]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc529_phy_pc_w))
                begin
                    if(good[long_cpuid529/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid529 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid529/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid529])
        end // if (done[529])

        if (done[530]) begin
            timeout[long_cpuid530] = 0;
            //check_bad_trap(spc530_phy_pc_w, 530, long_cpuid530);
            if(active_thread[long_cpuid530])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc530_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid530/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 530 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid530]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc530_phy_pc_w))
                begin
                    if(good[long_cpuid530/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid530 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid530/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid530])
        end // if (done[530])

        if (done[531]) begin
            timeout[long_cpuid531] = 0;
            //check_bad_trap(spc531_phy_pc_w, 531, long_cpuid531);
            if(active_thread[long_cpuid531])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc531_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid531/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 531 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid531]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc531_phy_pc_w))
                begin
                    if(good[long_cpuid531/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid531 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid531/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid531])
        end // if (done[531])

        if (done[532]) begin
            timeout[long_cpuid532] = 0;
            //check_bad_trap(spc532_phy_pc_w, 532, long_cpuid532);
            if(active_thread[long_cpuid532])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc532_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid532/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 532 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid532]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc532_phy_pc_w))
                begin
                    if(good[long_cpuid532/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid532 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid532/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid532])
        end // if (done[532])

        if (done[533]) begin
            timeout[long_cpuid533] = 0;
            //check_bad_trap(spc533_phy_pc_w, 533, long_cpuid533);
            if(active_thread[long_cpuid533])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc533_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid533/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 533 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid533]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc533_phy_pc_w))
                begin
                    if(good[long_cpuid533/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid533 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid533/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid533])
        end // if (done[533])

        if (done[534]) begin
            timeout[long_cpuid534] = 0;
            //check_bad_trap(spc534_phy_pc_w, 534, long_cpuid534);
            if(active_thread[long_cpuid534])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc534_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid534/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 534 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid534]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc534_phy_pc_w))
                begin
                    if(good[long_cpuid534/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid534 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid534/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid534])
        end // if (done[534])

        if (done[535]) begin
            timeout[long_cpuid535] = 0;
            //check_bad_trap(spc535_phy_pc_w, 535, long_cpuid535);
            if(active_thread[long_cpuid535])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc535_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid535/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 535 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid535]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc535_phy_pc_w))
                begin
                    if(good[long_cpuid535/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid535 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid535/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid535])
        end // if (done[535])

        if (done[536]) begin
            timeout[long_cpuid536] = 0;
            //check_bad_trap(spc536_phy_pc_w, 536, long_cpuid536);
            if(active_thread[long_cpuid536])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc536_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid536/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 536 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid536]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc536_phy_pc_w))
                begin
                    if(good[long_cpuid536/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid536 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid536/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid536])
        end // if (done[536])

        if (done[537]) begin
            timeout[long_cpuid537] = 0;
            //check_bad_trap(spc537_phy_pc_w, 537, long_cpuid537);
            if(active_thread[long_cpuid537])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc537_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid537/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 537 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid537]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc537_phy_pc_w))
                begin
                    if(good[long_cpuid537/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid537 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid537/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid537])
        end // if (done[537])

        if (done[538]) begin
            timeout[long_cpuid538] = 0;
            //check_bad_trap(spc538_phy_pc_w, 538, long_cpuid538);
            if(active_thread[long_cpuid538])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc538_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid538/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 538 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid538]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc538_phy_pc_w))
                begin
                    if(good[long_cpuid538/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid538 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid538/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid538])
        end // if (done[538])

        if (done[539]) begin
            timeout[long_cpuid539] = 0;
            //check_bad_trap(spc539_phy_pc_w, 539, long_cpuid539);
            if(active_thread[long_cpuid539])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc539_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid539/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 539 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid539]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc539_phy_pc_w))
                begin
                    if(good[long_cpuid539/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid539 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid539/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid539])
        end // if (done[539])

        if (done[540]) begin
            timeout[long_cpuid540] = 0;
            //check_bad_trap(spc540_phy_pc_w, 540, long_cpuid540);
            if(active_thread[long_cpuid540])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc540_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid540/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 540 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid540]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc540_phy_pc_w))
                begin
                    if(good[long_cpuid540/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid540 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid540/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid540])
        end // if (done[540])

        if (done[541]) begin
            timeout[long_cpuid541] = 0;
            //check_bad_trap(spc541_phy_pc_w, 541, long_cpuid541);
            if(active_thread[long_cpuid541])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc541_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid541/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 541 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid541]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc541_phy_pc_w))
                begin
                    if(good[long_cpuid541/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid541 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid541/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid541])
        end // if (done[541])

        if (done[542]) begin
            timeout[long_cpuid542] = 0;
            //check_bad_trap(spc542_phy_pc_w, 542, long_cpuid542);
            if(active_thread[long_cpuid542])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc542_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid542/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 542 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid542]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc542_phy_pc_w))
                begin
                    if(good[long_cpuid542/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid542 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid542/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid542])
        end // if (done[542])

        if (done[543]) begin
            timeout[long_cpuid543] = 0;
            //check_bad_trap(spc543_phy_pc_w, 543, long_cpuid543);
            if(active_thread[long_cpuid543])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc543_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid543/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 543 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid543]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc543_phy_pc_w))
                begin
                    if(good[long_cpuid543/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid543 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid543/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid543])
        end // if (done[543])

        if (done[544]) begin
            timeout[long_cpuid544] = 0;
            //check_bad_trap(spc544_phy_pc_w, 544, long_cpuid544);
            if(active_thread[long_cpuid544])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc544_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid544/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 544 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid544]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc544_phy_pc_w))
                begin
                    if(good[long_cpuid544/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid544 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid544/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid544])
        end // if (done[544])

        if (done[545]) begin
            timeout[long_cpuid545] = 0;
            //check_bad_trap(spc545_phy_pc_w, 545, long_cpuid545);
            if(active_thread[long_cpuid545])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc545_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid545/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 545 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid545]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc545_phy_pc_w))
                begin
                    if(good[long_cpuid545/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid545 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid545/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid545])
        end // if (done[545])

        if (done[546]) begin
            timeout[long_cpuid546] = 0;
            //check_bad_trap(spc546_phy_pc_w, 546, long_cpuid546);
            if(active_thread[long_cpuid546])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc546_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid546/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 546 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid546]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc546_phy_pc_w))
                begin
                    if(good[long_cpuid546/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid546 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid546/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid546])
        end // if (done[546])

        if (done[547]) begin
            timeout[long_cpuid547] = 0;
            //check_bad_trap(spc547_phy_pc_w, 547, long_cpuid547);
            if(active_thread[long_cpuid547])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc547_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid547/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 547 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid547]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc547_phy_pc_w))
                begin
                    if(good[long_cpuid547/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid547 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid547/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid547])
        end // if (done[547])

        if (done[548]) begin
            timeout[long_cpuid548] = 0;
            //check_bad_trap(spc548_phy_pc_w, 548, long_cpuid548);
            if(active_thread[long_cpuid548])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc548_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid548/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 548 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid548]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc548_phy_pc_w))
                begin
                    if(good[long_cpuid548/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid548 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid548/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid548])
        end // if (done[548])

        if (done[549]) begin
            timeout[long_cpuid549] = 0;
            //check_bad_trap(spc549_phy_pc_w, 549, long_cpuid549);
            if(active_thread[long_cpuid549])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc549_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid549/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 549 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid549]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc549_phy_pc_w))
                begin
                    if(good[long_cpuid549/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid549 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid549/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid549])
        end // if (done[549])

        if (done[550]) begin
            timeout[long_cpuid550] = 0;
            //check_bad_trap(spc550_phy_pc_w, 550, long_cpuid550);
            if(active_thread[long_cpuid550])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc550_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid550/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 550 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid550]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc550_phy_pc_w))
                begin
                    if(good[long_cpuid550/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid550 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid550/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid550])
        end // if (done[550])

        if (done[551]) begin
            timeout[long_cpuid551] = 0;
            //check_bad_trap(spc551_phy_pc_w, 551, long_cpuid551);
            if(active_thread[long_cpuid551])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc551_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid551/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 551 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid551]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc551_phy_pc_w))
                begin
                    if(good[long_cpuid551/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid551 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid551/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid551])
        end // if (done[551])

        if (done[552]) begin
            timeout[long_cpuid552] = 0;
            //check_bad_trap(spc552_phy_pc_w, 552, long_cpuid552);
            if(active_thread[long_cpuid552])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc552_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid552/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 552 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid552]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc552_phy_pc_w))
                begin
                    if(good[long_cpuid552/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid552 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid552/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid552])
        end // if (done[552])

        if (done[553]) begin
            timeout[long_cpuid553] = 0;
            //check_bad_trap(spc553_phy_pc_w, 553, long_cpuid553);
            if(active_thread[long_cpuid553])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc553_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid553/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 553 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid553]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc553_phy_pc_w))
                begin
                    if(good[long_cpuid553/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid553 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid553/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid553])
        end // if (done[553])

        if (done[554]) begin
            timeout[long_cpuid554] = 0;
            //check_bad_trap(spc554_phy_pc_w, 554, long_cpuid554);
            if(active_thread[long_cpuid554])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc554_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid554/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 554 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid554]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc554_phy_pc_w))
                begin
                    if(good[long_cpuid554/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid554 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid554/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid554])
        end // if (done[554])

        if (done[555]) begin
            timeout[long_cpuid555] = 0;
            //check_bad_trap(spc555_phy_pc_w, 555, long_cpuid555);
            if(active_thread[long_cpuid555])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc555_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid555/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 555 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid555]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc555_phy_pc_w))
                begin
                    if(good[long_cpuid555/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid555 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid555/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid555])
        end // if (done[555])

        if (done[556]) begin
            timeout[long_cpuid556] = 0;
            //check_bad_trap(spc556_phy_pc_w, 556, long_cpuid556);
            if(active_thread[long_cpuid556])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc556_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid556/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 556 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid556]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc556_phy_pc_w))
                begin
                    if(good[long_cpuid556/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid556 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid556/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid556])
        end // if (done[556])

        if (done[557]) begin
            timeout[long_cpuid557] = 0;
            //check_bad_trap(spc557_phy_pc_w, 557, long_cpuid557);
            if(active_thread[long_cpuid557])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc557_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid557/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 557 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid557]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc557_phy_pc_w))
                begin
                    if(good[long_cpuid557/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid557 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid557/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid557])
        end // if (done[557])

        if (done[558]) begin
            timeout[long_cpuid558] = 0;
            //check_bad_trap(spc558_phy_pc_w, 558, long_cpuid558);
            if(active_thread[long_cpuid558])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc558_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid558/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 558 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid558]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc558_phy_pc_w))
                begin
                    if(good[long_cpuid558/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid558 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid558/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid558])
        end // if (done[558])

        if (done[559]) begin
            timeout[long_cpuid559] = 0;
            //check_bad_trap(spc559_phy_pc_w, 559, long_cpuid559);
            if(active_thread[long_cpuid559])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc559_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid559/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 559 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid559]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc559_phy_pc_w))
                begin
                    if(good[long_cpuid559/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid559 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid559/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid559])
        end // if (done[559])

        if (done[560]) begin
            timeout[long_cpuid560] = 0;
            //check_bad_trap(spc560_phy_pc_w, 560, long_cpuid560);
            if(active_thread[long_cpuid560])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc560_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid560/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 560 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid560]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc560_phy_pc_w))
                begin
                    if(good[long_cpuid560/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid560 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid560/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid560])
        end // if (done[560])

        if (done[561]) begin
            timeout[long_cpuid561] = 0;
            //check_bad_trap(spc561_phy_pc_w, 561, long_cpuid561);
            if(active_thread[long_cpuid561])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc561_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid561/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 561 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid561]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc561_phy_pc_w))
                begin
                    if(good[long_cpuid561/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid561 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid561/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid561])
        end // if (done[561])

        if (done[562]) begin
            timeout[long_cpuid562] = 0;
            //check_bad_trap(spc562_phy_pc_w, 562, long_cpuid562);
            if(active_thread[long_cpuid562])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc562_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid562/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 562 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid562]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc562_phy_pc_w))
                begin
                    if(good[long_cpuid562/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid562 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid562/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid562])
        end // if (done[562])

        if (done[563]) begin
            timeout[long_cpuid563] = 0;
            //check_bad_trap(spc563_phy_pc_w, 563, long_cpuid563);
            if(active_thread[long_cpuid563])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc563_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid563/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 563 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid563]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc563_phy_pc_w))
                begin
                    if(good[long_cpuid563/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid563 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid563/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid563])
        end // if (done[563])

        if (done[564]) begin
            timeout[long_cpuid564] = 0;
            //check_bad_trap(spc564_phy_pc_w, 564, long_cpuid564);
            if(active_thread[long_cpuid564])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc564_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid564/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 564 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid564]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc564_phy_pc_w))
                begin
                    if(good[long_cpuid564/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid564 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid564/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid564])
        end // if (done[564])

        if (done[565]) begin
            timeout[long_cpuid565] = 0;
            //check_bad_trap(spc565_phy_pc_w, 565, long_cpuid565);
            if(active_thread[long_cpuid565])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc565_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid565/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 565 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid565]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc565_phy_pc_w))
                begin
                    if(good[long_cpuid565/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid565 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid565/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid565])
        end // if (done[565])

        if (done[566]) begin
            timeout[long_cpuid566] = 0;
            //check_bad_trap(spc566_phy_pc_w, 566, long_cpuid566);
            if(active_thread[long_cpuid566])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc566_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid566/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 566 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid566]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc566_phy_pc_w))
                begin
                    if(good[long_cpuid566/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid566 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid566/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid566])
        end // if (done[566])

        if (done[567]) begin
            timeout[long_cpuid567] = 0;
            //check_bad_trap(spc567_phy_pc_w, 567, long_cpuid567);
            if(active_thread[long_cpuid567])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc567_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid567/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 567 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid567]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc567_phy_pc_w))
                begin
                    if(good[long_cpuid567/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid567 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid567/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid567])
        end // if (done[567])

        if (done[568]) begin
            timeout[long_cpuid568] = 0;
            //check_bad_trap(spc568_phy_pc_w, 568, long_cpuid568);
            if(active_thread[long_cpuid568])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc568_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid568/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 568 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid568]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc568_phy_pc_w))
                begin
                    if(good[long_cpuid568/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid568 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid568/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid568])
        end // if (done[568])

        if (done[569]) begin
            timeout[long_cpuid569] = 0;
            //check_bad_trap(spc569_phy_pc_w, 569, long_cpuid569);
            if(active_thread[long_cpuid569])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc569_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid569/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 569 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid569]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc569_phy_pc_w))
                begin
                    if(good[long_cpuid569/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid569 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid569/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid569])
        end // if (done[569])

        if (done[570]) begin
            timeout[long_cpuid570] = 0;
            //check_bad_trap(spc570_phy_pc_w, 570, long_cpuid570);
            if(active_thread[long_cpuid570])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc570_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid570/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 570 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid570]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc570_phy_pc_w))
                begin
                    if(good[long_cpuid570/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid570 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid570/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid570])
        end // if (done[570])

        if (done[571]) begin
            timeout[long_cpuid571] = 0;
            //check_bad_trap(spc571_phy_pc_w, 571, long_cpuid571);
            if(active_thread[long_cpuid571])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc571_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid571/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 571 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid571]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc571_phy_pc_w))
                begin
                    if(good[long_cpuid571/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid571 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid571/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid571])
        end // if (done[571])

        if (done[572]) begin
            timeout[long_cpuid572] = 0;
            //check_bad_trap(spc572_phy_pc_w, 572, long_cpuid572);
            if(active_thread[long_cpuid572])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc572_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid572/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 572 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid572]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc572_phy_pc_w))
                begin
                    if(good[long_cpuid572/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid572 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid572/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid572])
        end // if (done[572])

        if (done[573]) begin
            timeout[long_cpuid573] = 0;
            //check_bad_trap(spc573_phy_pc_w, 573, long_cpuid573);
            if(active_thread[long_cpuid573])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc573_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid573/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 573 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid573]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc573_phy_pc_w))
                begin
                    if(good[long_cpuid573/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid573 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid573/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid573])
        end // if (done[573])

        if (done[574]) begin
            timeout[long_cpuid574] = 0;
            //check_bad_trap(spc574_phy_pc_w, 574, long_cpuid574);
            if(active_thread[long_cpuid574])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc574_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid574/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 574 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid574]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc574_phy_pc_w))
                begin
                    if(good[long_cpuid574/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid574 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid574/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid574])
        end // if (done[574])

        if (done[575]) begin
            timeout[long_cpuid575] = 0;
            //check_bad_trap(spc575_phy_pc_w, 575, long_cpuid575);
            if(active_thread[long_cpuid575])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc575_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid575/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 575 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid575]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc575_phy_pc_w))
                begin
                    if(good[long_cpuid575/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid575 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid575/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid575])
        end // if (done[575])

        if (done[576]) begin
            timeout[long_cpuid576] = 0;
            //check_bad_trap(spc576_phy_pc_w, 576, long_cpuid576);
            if(active_thread[long_cpuid576])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc576_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid576/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 576 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid576]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc576_phy_pc_w))
                begin
                    if(good[long_cpuid576/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid576 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid576/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid576])
        end // if (done[576])

        if (done[577]) begin
            timeout[long_cpuid577] = 0;
            //check_bad_trap(spc577_phy_pc_w, 577, long_cpuid577);
            if(active_thread[long_cpuid577])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc577_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid577/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 577 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid577]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc577_phy_pc_w))
                begin
                    if(good[long_cpuid577/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid577 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid577/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid577])
        end // if (done[577])

        if (done[578]) begin
            timeout[long_cpuid578] = 0;
            //check_bad_trap(spc578_phy_pc_w, 578, long_cpuid578);
            if(active_thread[long_cpuid578])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc578_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid578/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 578 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid578]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc578_phy_pc_w))
                begin
                    if(good[long_cpuid578/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid578 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid578/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid578])
        end // if (done[578])

        if (done[579]) begin
            timeout[long_cpuid579] = 0;
            //check_bad_trap(spc579_phy_pc_w, 579, long_cpuid579);
            if(active_thread[long_cpuid579])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc579_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid579/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 579 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid579]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc579_phy_pc_w))
                begin
                    if(good[long_cpuid579/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid579 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid579/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid579])
        end // if (done[579])

        if (done[580]) begin
            timeout[long_cpuid580] = 0;
            //check_bad_trap(spc580_phy_pc_w, 580, long_cpuid580);
            if(active_thread[long_cpuid580])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc580_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid580/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 580 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid580]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc580_phy_pc_w))
                begin
                    if(good[long_cpuid580/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid580 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid580/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid580])
        end // if (done[580])

        if (done[581]) begin
            timeout[long_cpuid581] = 0;
            //check_bad_trap(spc581_phy_pc_w, 581, long_cpuid581);
            if(active_thread[long_cpuid581])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc581_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid581/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 581 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid581]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc581_phy_pc_w))
                begin
                    if(good[long_cpuid581/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid581 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid581/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid581])
        end // if (done[581])

        if (done[582]) begin
            timeout[long_cpuid582] = 0;
            //check_bad_trap(spc582_phy_pc_w, 582, long_cpuid582);
            if(active_thread[long_cpuid582])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc582_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid582/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 582 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid582]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc582_phy_pc_w))
                begin
                    if(good[long_cpuid582/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid582 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid582/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid582])
        end // if (done[582])

        if (done[583]) begin
            timeout[long_cpuid583] = 0;
            //check_bad_trap(spc583_phy_pc_w, 583, long_cpuid583);
            if(active_thread[long_cpuid583])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc583_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid583/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 583 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid583]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc583_phy_pc_w))
                begin
                    if(good[long_cpuid583/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid583 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid583/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid583])
        end // if (done[583])

        if (done[584]) begin
            timeout[long_cpuid584] = 0;
            //check_bad_trap(spc584_phy_pc_w, 584, long_cpuid584);
            if(active_thread[long_cpuid584])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc584_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid584/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 584 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid584]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc584_phy_pc_w))
                begin
                    if(good[long_cpuid584/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid584 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid584/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid584])
        end // if (done[584])

        if (done[585]) begin
            timeout[long_cpuid585] = 0;
            //check_bad_trap(spc585_phy_pc_w, 585, long_cpuid585);
            if(active_thread[long_cpuid585])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc585_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid585/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 585 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid585]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc585_phy_pc_w))
                begin
                    if(good[long_cpuid585/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid585 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid585/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid585])
        end // if (done[585])

        if (done[586]) begin
            timeout[long_cpuid586] = 0;
            //check_bad_trap(spc586_phy_pc_w, 586, long_cpuid586);
            if(active_thread[long_cpuid586])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc586_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid586/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 586 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid586]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc586_phy_pc_w))
                begin
                    if(good[long_cpuid586/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid586 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid586/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid586])
        end // if (done[586])

        if (done[587]) begin
            timeout[long_cpuid587] = 0;
            //check_bad_trap(spc587_phy_pc_w, 587, long_cpuid587);
            if(active_thread[long_cpuid587])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc587_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid587/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 587 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid587]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc587_phy_pc_w))
                begin
                    if(good[long_cpuid587/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid587 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid587/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid587])
        end // if (done[587])

        if (done[588]) begin
            timeout[long_cpuid588] = 0;
            //check_bad_trap(spc588_phy_pc_w, 588, long_cpuid588);
            if(active_thread[long_cpuid588])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc588_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid588/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 588 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid588]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc588_phy_pc_w))
                begin
                    if(good[long_cpuid588/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid588 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid588/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid588])
        end // if (done[588])

        if (done[589]) begin
            timeout[long_cpuid589] = 0;
            //check_bad_trap(spc589_phy_pc_w, 589, long_cpuid589);
            if(active_thread[long_cpuid589])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc589_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid589/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 589 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid589]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc589_phy_pc_w))
                begin
                    if(good[long_cpuid589/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid589 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid589/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid589])
        end // if (done[589])

        if (done[590]) begin
            timeout[long_cpuid590] = 0;
            //check_bad_trap(spc590_phy_pc_w, 590, long_cpuid590);
            if(active_thread[long_cpuid590])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc590_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid590/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 590 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid590]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc590_phy_pc_w))
                begin
                    if(good[long_cpuid590/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid590 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid590/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid590])
        end // if (done[590])

        if (done[591]) begin
            timeout[long_cpuid591] = 0;
            //check_bad_trap(spc591_phy_pc_w, 591, long_cpuid591);
            if(active_thread[long_cpuid591])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc591_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid591/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 591 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid591]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc591_phy_pc_w))
                begin
                    if(good[long_cpuid591/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid591 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid591/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid591])
        end // if (done[591])

        if (done[592]) begin
            timeout[long_cpuid592] = 0;
            //check_bad_trap(spc592_phy_pc_w, 592, long_cpuid592);
            if(active_thread[long_cpuid592])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc592_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid592/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 592 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid592]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc592_phy_pc_w))
                begin
                    if(good[long_cpuid592/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid592 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid592/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid592])
        end // if (done[592])

        if (done[593]) begin
            timeout[long_cpuid593] = 0;
            //check_bad_trap(spc593_phy_pc_w, 593, long_cpuid593);
            if(active_thread[long_cpuid593])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc593_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid593/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 593 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid593]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc593_phy_pc_w))
                begin
                    if(good[long_cpuid593/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid593 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid593/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid593])
        end // if (done[593])

        if (done[594]) begin
            timeout[long_cpuid594] = 0;
            //check_bad_trap(spc594_phy_pc_w, 594, long_cpuid594);
            if(active_thread[long_cpuid594])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc594_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid594/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 594 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid594]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc594_phy_pc_w))
                begin
                    if(good[long_cpuid594/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid594 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid594/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid594])
        end // if (done[594])

        if (done[595]) begin
            timeout[long_cpuid595] = 0;
            //check_bad_trap(spc595_phy_pc_w, 595, long_cpuid595);
            if(active_thread[long_cpuid595])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc595_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid595/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 595 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid595]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc595_phy_pc_w))
                begin
                    if(good[long_cpuid595/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid595 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid595/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid595])
        end // if (done[595])

        if (done[596]) begin
            timeout[long_cpuid596] = 0;
            //check_bad_trap(spc596_phy_pc_w, 596, long_cpuid596);
            if(active_thread[long_cpuid596])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc596_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid596/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 596 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid596]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc596_phy_pc_w))
                begin
                    if(good[long_cpuid596/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid596 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid596/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid596])
        end // if (done[596])

        if (done[597]) begin
            timeout[long_cpuid597] = 0;
            //check_bad_trap(spc597_phy_pc_w, 597, long_cpuid597);
            if(active_thread[long_cpuid597])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc597_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid597/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 597 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid597]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc597_phy_pc_w))
                begin
                    if(good[long_cpuid597/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid597 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid597/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid597])
        end // if (done[597])

        if (done[598]) begin
            timeout[long_cpuid598] = 0;
            //check_bad_trap(spc598_phy_pc_w, 598, long_cpuid598);
            if(active_thread[long_cpuid598])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc598_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid598/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 598 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid598]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc598_phy_pc_w))
                begin
                    if(good[long_cpuid598/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid598 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid598/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid598])
        end // if (done[598])

        if (done[599]) begin
            timeout[long_cpuid599] = 0;
            //check_bad_trap(spc599_phy_pc_w, 599, long_cpuid599);
            if(active_thread[long_cpuid599])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc599_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid599/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 599 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid599]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc599_phy_pc_w))
                begin
                    if(good[long_cpuid599/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid599 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid599/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid599])
        end // if (done[599])

        if (done[600]) begin
            timeout[long_cpuid600] = 0;
            //check_bad_trap(spc600_phy_pc_w, 600, long_cpuid600);
            if(active_thread[long_cpuid600])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc600_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid600/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 600 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid600]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc600_phy_pc_w))
                begin
                    if(good[long_cpuid600/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid600 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid600/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid600])
        end // if (done[600])

        if (done[601]) begin
            timeout[long_cpuid601] = 0;
            //check_bad_trap(spc601_phy_pc_w, 601, long_cpuid601);
            if(active_thread[long_cpuid601])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc601_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid601/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 601 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid601]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc601_phy_pc_w))
                begin
                    if(good[long_cpuid601/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid601 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid601/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid601])
        end // if (done[601])

        if (done[602]) begin
            timeout[long_cpuid602] = 0;
            //check_bad_trap(spc602_phy_pc_w, 602, long_cpuid602);
            if(active_thread[long_cpuid602])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc602_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid602/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 602 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid602]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc602_phy_pc_w))
                begin
                    if(good[long_cpuid602/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid602 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid602/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid602])
        end // if (done[602])

        if (done[603]) begin
            timeout[long_cpuid603] = 0;
            //check_bad_trap(spc603_phy_pc_w, 603, long_cpuid603);
            if(active_thread[long_cpuid603])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc603_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid603/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 603 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid603]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc603_phy_pc_w))
                begin
                    if(good[long_cpuid603/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid603 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid603/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid603])
        end // if (done[603])

        if (done[604]) begin
            timeout[long_cpuid604] = 0;
            //check_bad_trap(spc604_phy_pc_w, 604, long_cpuid604);
            if(active_thread[long_cpuid604])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc604_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid604/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 604 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid604]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc604_phy_pc_w))
                begin
                    if(good[long_cpuid604/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid604 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid604/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid604])
        end // if (done[604])

        if (done[605]) begin
            timeout[long_cpuid605] = 0;
            //check_bad_trap(spc605_phy_pc_w, 605, long_cpuid605);
            if(active_thread[long_cpuid605])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc605_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid605/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 605 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid605]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc605_phy_pc_w))
                begin
                    if(good[long_cpuid605/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid605 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid605/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid605])
        end // if (done[605])

        if (done[606]) begin
            timeout[long_cpuid606] = 0;
            //check_bad_trap(spc606_phy_pc_w, 606, long_cpuid606);
            if(active_thread[long_cpuid606])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc606_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid606/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 606 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid606]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc606_phy_pc_w))
                begin
                    if(good[long_cpuid606/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid606 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid606/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid606])
        end // if (done[606])

        if (done[607]) begin
            timeout[long_cpuid607] = 0;
            //check_bad_trap(spc607_phy_pc_w, 607, long_cpuid607);
            if(active_thread[long_cpuid607])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc607_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid607/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 607 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid607]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc607_phy_pc_w))
                begin
                    if(good[long_cpuid607/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid607 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid607/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid607])
        end // if (done[607])

        if (done[608]) begin
            timeout[long_cpuid608] = 0;
            //check_bad_trap(spc608_phy_pc_w, 608, long_cpuid608);
            if(active_thread[long_cpuid608])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc608_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid608/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 608 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid608]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc608_phy_pc_w))
                begin
                    if(good[long_cpuid608/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid608 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid608/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid608])
        end // if (done[608])

        if (done[609]) begin
            timeout[long_cpuid609] = 0;
            //check_bad_trap(spc609_phy_pc_w, 609, long_cpuid609);
            if(active_thread[long_cpuid609])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc609_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid609/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 609 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid609]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc609_phy_pc_w))
                begin
                    if(good[long_cpuid609/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid609 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid609/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid609])
        end // if (done[609])

        if (done[610]) begin
            timeout[long_cpuid610] = 0;
            //check_bad_trap(spc610_phy_pc_w, 610, long_cpuid610);
            if(active_thread[long_cpuid610])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc610_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid610/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 610 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid610]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc610_phy_pc_w))
                begin
                    if(good[long_cpuid610/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid610 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid610/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid610])
        end // if (done[610])

        if (done[611]) begin
            timeout[long_cpuid611] = 0;
            //check_bad_trap(spc611_phy_pc_w, 611, long_cpuid611);
            if(active_thread[long_cpuid611])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc611_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid611/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 611 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid611]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc611_phy_pc_w))
                begin
                    if(good[long_cpuid611/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid611 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid611/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid611])
        end // if (done[611])

        if (done[612]) begin
            timeout[long_cpuid612] = 0;
            //check_bad_trap(spc612_phy_pc_w, 612, long_cpuid612);
            if(active_thread[long_cpuid612])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc612_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid612/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 612 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid612]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc612_phy_pc_w))
                begin
                    if(good[long_cpuid612/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid612 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid612/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid612])
        end // if (done[612])

        if (done[613]) begin
            timeout[long_cpuid613] = 0;
            //check_bad_trap(spc613_phy_pc_w, 613, long_cpuid613);
            if(active_thread[long_cpuid613])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc613_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid613/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 613 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid613]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc613_phy_pc_w))
                begin
                    if(good[long_cpuid613/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid613 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid613/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid613])
        end // if (done[613])

        if (done[614]) begin
            timeout[long_cpuid614] = 0;
            //check_bad_trap(spc614_phy_pc_w, 614, long_cpuid614);
            if(active_thread[long_cpuid614])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc614_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid614/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 614 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid614]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc614_phy_pc_w))
                begin
                    if(good[long_cpuid614/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid614 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid614/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid614])
        end // if (done[614])

        if (done[615]) begin
            timeout[long_cpuid615] = 0;
            //check_bad_trap(spc615_phy_pc_w, 615, long_cpuid615);
            if(active_thread[long_cpuid615])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc615_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid615/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 615 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid615]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc615_phy_pc_w))
                begin
                    if(good[long_cpuid615/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid615 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid615/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid615])
        end // if (done[615])

        if (done[616]) begin
            timeout[long_cpuid616] = 0;
            //check_bad_trap(spc616_phy_pc_w, 616, long_cpuid616);
            if(active_thread[long_cpuid616])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc616_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid616/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 616 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid616]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc616_phy_pc_w))
                begin
                    if(good[long_cpuid616/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid616 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid616/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid616])
        end // if (done[616])

        if (done[617]) begin
            timeout[long_cpuid617] = 0;
            //check_bad_trap(spc617_phy_pc_w, 617, long_cpuid617);
            if(active_thread[long_cpuid617])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc617_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid617/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 617 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid617]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc617_phy_pc_w))
                begin
                    if(good[long_cpuid617/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid617 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid617/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid617])
        end // if (done[617])

        if (done[618]) begin
            timeout[long_cpuid618] = 0;
            //check_bad_trap(spc618_phy_pc_w, 618, long_cpuid618);
            if(active_thread[long_cpuid618])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc618_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid618/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 618 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid618]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc618_phy_pc_w))
                begin
                    if(good[long_cpuid618/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid618 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid618/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid618])
        end // if (done[618])

        if (done[619]) begin
            timeout[long_cpuid619] = 0;
            //check_bad_trap(spc619_phy_pc_w, 619, long_cpuid619);
            if(active_thread[long_cpuid619])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc619_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid619/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 619 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid619]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc619_phy_pc_w))
                begin
                    if(good[long_cpuid619/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid619 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid619/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid619])
        end // if (done[619])

        if (done[620]) begin
            timeout[long_cpuid620] = 0;
            //check_bad_trap(spc620_phy_pc_w, 620, long_cpuid620);
            if(active_thread[long_cpuid620])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc620_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid620/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 620 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid620]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc620_phy_pc_w))
                begin
                    if(good[long_cpuid620/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid620 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid620/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid620])
        end // if (done[620])

        if (done[621]) begin
            timeout[long_cpuid621] = 0;
            //check_bad_trap(spc621_phy_pc_w, 621, long_cpuid621);
            if(active_thread[long_cpuid621])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc621_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid621/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 621 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid621]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc621_phy_pc_w))
                begin
                    if(good[long_cpuid621/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid621 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid621/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid621])
        end // if (done[621])

        if (done[622]) begin
            timeout[long_cpuid622] = 0;
            //check_bad_trap(spc622_phy_pc_w, 622, long_cpuid622);
            if(active_thread[long_cpuid622])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc622_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid622/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 622 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid622]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc622_phy_pc_w))
                begin
                    if(good[long_cpuid622/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid622 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid622/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid622])
        end // if (done[622])

        if (done[623]) begin
            timeout[long_cpuid623] = 0;
            //check_bad_trap(spc623_phy_pc_w, 623, long_cpuid623);
            if(active_thread[long_cpuid623])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc623_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid623/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 623 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid623]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc623_phy_pc_w))
                begin
                    if(good[long_cpuid623/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid623 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid623/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid623])
        end // if (done[623])

        if (done[624]) begin
            timeout[long_cpuid624] = 0;
            //check_bad_trap(spc624_phy_pc_w, 624, long_cpuid624);
            if(active_thread[long_cpuid624])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc624_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid624/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 624 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid624]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc624_phy_pc_w))
                begin
                    if(good[long_cpuid624/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid624 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid624/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid624])
        end // if (done[624])

        if (done[625]) begin
            timeout[long_cpuid625] = 0;
            //check_bad_trap(spc625_phy_pc_w, 625, long_cpuid625);
            if(active_thread[long_cpuid625])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc625_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid625/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 625 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid625]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc625_phy_pc_w))
                begin
                    if(good[long_cpuid625/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid625 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid625/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid625])
        end // if (done[625])

        if (done[626]) begin
            timeout[long_cpuid626] = 0;
            //check_bad_trap(spc626_phy_pc_w, 626, long_cpuid626);
            if(active_thread[long_cpuid626])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc626_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid626/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 626 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid626]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc626_phy_pc_w))
                begin
                    if(good[long_cpuid626/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid626 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid626/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid626])
        end // if (done[626])

        if (done[627]) begin
            timeout[long_cpuid627] = 0;
            //check_bad_trap(spc627_phy_pc_w, 627, long_cpuid627);
            if(active_thread[long_cpuid627])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc627_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid627/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 627 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid627]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc627_phy_pc_w))
                begin
                    if(good[long_cpuid627/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid627 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid627/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid627])
        end // if (done[627])

        if (done[628]) begin
            timeout[long_cpuid628] = 0;
            //check_bad_trap(spc628_phy_pc_w, 628, long_cpuid628);
            if(active_thread[long_cpuid628])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc628_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid628/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 628 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid628]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc628_phy_pc_w))
                begin
                    if(good[long_cpuid628/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid628 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid628/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid628])
        end // if (done[628])

        if (done[629]) begin
            timeout[long_cpuid629] = 0;
            //check_bad_trap(spc629_phy_pc_w, 629, long_cpuid629);
            if(active_thread[long_cpuid629])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc629_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid629/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 629 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid629]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc629_phy_pc_w))
                begin
                    if(good[long_cpuid629/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid629 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid629/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid629])
        end // if (done[629])

        if (done[630]) begin
            timeout[long_cpuid630] = 0;
            //check_bad_trap(spc630_phy_pc_w, 630, long_cpuid630);
            if(active_thread[long_cpuid630])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc630_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid630/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 630 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid630]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc630_phy_pc_w))
                begin
                    if(good[long_cpuid630/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid630 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid630/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid630])
        end // if (done[630])

        if (done[631]) begin
            timeout[long_cpuid631] = 0;
            //check_bad_trap(spc631_phy_pc_w, 631, long_cpuid631);
            if(active_thread[long_cpuid631])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc631_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid631/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 631 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid631]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc631_phy_pc_w))
                begin
                    if(good[long_cpuid631/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid631 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid631/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid631])
        end // if (done[631])

        if (done[632]) begin
            timeout[long_cpuid632] = 0;
            //check_bad_trap(spc632_phy_pc_w, 632, long_cpuid632);
            if(active_thread[long_cpuid632])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc632_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid632/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 632 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid632]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc632_phy_pc_w))
                begin
                    if(good[long_cpuid632/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid632 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid632/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid632])
        end // if (done[632])

        if (done[633]) begin
            timeout[long_cpuid633] = 0;
            //check_bad_trap(spc633_phy_pc_w, 633, long_cpuid633);
            if(active_thread[long_cpuid633])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc633_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid633/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 633 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid633]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc633_phy_pc_w))
                begin
                    if(good[long_cpuid633/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid633 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid633/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid633])
        end // if (done[633])

        if (done[634]) begin
            timeout[long_cpuid634] = 0;
            //check_bad_trap(spc634_phy_pc_w, 634, long_cpuid634);
            if(active_thread[long_cpuid634])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc634_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid634/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 634 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid634]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc634_phy_pc_w))
                begin
                    if(good[long_cpuid634/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid634 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid634/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid634])
        end // if (done[634])

        if (done[635]) begin
            timeout[long_cpuid635] = 0;
            //check_bad_trap(spc635_phy_pc_w, 635, long_cpuid635);
            if(active_thread[long_cpuid635])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc635_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid635/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 635 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid635]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc635_phy_pc_w))
                begin
                    if(good[long_cpuid635/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid635 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid635/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid635])
        end // if (done[635])

        if (done[636]) begin
            timeout[long_cpuid636] = 0;
            //check_bad_trap(spc636_phy_pc_w, 636, long_cpuid636);
            if(active_thread[long_cpuid636])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc636_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid636/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 636 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid636]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc636_phy_pc_w))
                begin
                    if(good[long_cpuid636/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid636 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid636/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid636])
        end // if (done[636])

        if (done[637]) begin
            timeout[long_cpuid637] = 0;
            //check_bad_trap(spc637_phy_pc_w, 637, long_cpuid637);
            if(active_thread[long_cpuid637])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc637_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid637/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 637 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid637]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc637_phy_pc_w))
                begin
                    if(good[long_cpuid637/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid637 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid637/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid637])
        end // if (done[637])

        if (done[638]) begin
            timeout[long_cpuid638] = 0;
            //check_bad_trap(spc638_phy_pc_w, 638, long_cpuid638);
            if(active_thread[long_cpuid638])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc638_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid638/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 638 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid638]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc638_phy_pc_w))
                begin
                    if(good[long_cpuid638/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid638 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid638/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid638])
        end // if (done[638])

        if (done[639]) begin
            timeout[long_cpuid639] = 0;
            //check_bad_trap(spc639_phy_pc_w, 639, long_cpuid639);
            if(active_thread[long_cpuid639])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc639_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid639/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 639 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid639]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc639_phy_pc_w))
                begin
                    if(good[long_cpuid639/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid639 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid639/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid639])
        end // if (done[639])

        if (done[640]) begin
            timeout[long_cpuid640] = 0;
            //check_bad_trap(spc640_phy_pc_w, 640, long_cpuid640);
            if(active_thread[long_cpuid640])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc640_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid640/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 640 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid640]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc640_phy_pc_w))
                begin
                    if(good[long_cpuid640/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid640 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid640/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid640])
        end // if (done[640])

        if (done[641]) begin
            timeout[long_cpuid641] = 0;
            //check_bad_trap(spc641_phy_pc_w, 641, long_cpuid641);
            if(active_thread[long_cpuid641])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc641_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid641/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 641 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid641]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc641_phy_pc_w))
                begin
                    if(good[long_cpuid641/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid641 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid641/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid641])
        end // if (done[641])

        if (done[642]) begin
            timeout[long_cpuid642] = 0;
            //check_bad_trap(spc642_phy_pc_w, 642, long_cpuid642);
            if(active_thread[long_cpuid642])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc642_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid642/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 642 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid642]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc642_phy_pc_w))
                begin
                    if(good[long_cpuid642/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid642 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid642/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid642])
        end // if (done[642])

        if (done[643]) begin
            timeout[long_cpuid643] = 0;
            //check_bad_trap(spc643_phy_pc_w, 643, long_cpuid643);
            if(active_thread[long_cpuid643])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc643_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid643/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 643 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid643]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc643_phy_pc_w))
                begin
                    if(good[long_cpuid643/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid643 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid643/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid643])
        end // if (done[643])

        if (done[644]) begin
            timeout[long_cpuid644] = 0;
            //check_bad_trap(spc644_phy_pc_w, 644, long_cpuid644);
            if(active_thread[long_cpuid644])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc644_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid644/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 644 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid644]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc644_phy_pc_w))
                begin
                    if(good[long_cpuid644/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid644 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid644/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid644])
        end // if (done[644])

        if (done[645]) begin
            timeout[long_cpuid645] = 0;
            //check_bad_trap(spc645_phy_pc_w, 645, long_cpuid645);
            if(active_thread[long_cpuid645])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc645_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid645/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 645 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid645]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc645_phy_pc_w))
                begin
                    if(good[long_cpuid645/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid645 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid645/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid645])
        end // if (done[645])

        if (done[646]) begin
            timeout[long_cpuid646] = 0;
            //check_bad_trap(spc646_phy_pc_w, 646, long_cpuid646);
            if(active_thread[long_cpuid646])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc646_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid646/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 646 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid646]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc646_phy_pc_w))
                begin
                    if(good[long_cpuid646/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid646 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid646/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid646])
        end // if (done[646])

        if (done[647]) begin
            timeout[long_cpuid647] = 0;
            //check_bad_trap(spc647_phy_pc_w, 647, long_cpuid647);
            if(active_thread[long_cpuid647])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc647_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid647/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 647 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid647]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc647_phy_pc_w))
                begin
                    if(good[long_cpuid647/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid647 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid647/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid647])
        end // if (done[647])

        if (done[648]) begin
            timeout[long_cpuid648] = 0;
            //check_bad_trap(spc648_phy_pc_w, 648, long_cpuid648);
            if(active_thread[long_cpuid648])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc648_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid648/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 648 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid648]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc648_phy_pc_w))
                begin
                    if(good[long_cpuid648/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid648 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid648/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid648])
        end // if (done[648])

        if (done[649]) begin
            timeout[long_cpuid649] = 0;
            //check_bad_trap(spc649_phy_pc_w, 649, long_cpuid649);
            if(active_thread[long_cpuid649])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc649_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid649/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 649 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid649]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc649_phy_pc_w))
                begin
                    if(good[long_cpuid649/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid649 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid649/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid649])
        end // if (done[649])

        if (done[650]) begin
            timeout[long_cpuid650] = 0;
            //check_bad_trap(spc650_phy_pc_w, 650, long_cpuid650);
            if(active_thread[long_cpuid650])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc650_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid650/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 650 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid650]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc650_phy_pc_w))
                begin
                    if(good[long_cpuid650/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid650 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid650/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid650])
        end // if (done[650])

        if (done[651]) begin
            timeout[long_cpuid651] = 0;
            //check_bad_trap(spc651_phy_pc_w, 651, long_cpuid651);
            if(active_thread[long_cpuid651])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc651_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid651/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 651 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid651]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc651_phy_pc_w))
                begin
                    if(good[long_cpuid651/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid651 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid651/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid651])
        end // if (done[651])

        if (done[652]) begin
            timeout[long_cpuid652] = 0;
            //check_bad_trap(spc652_phy_pc_w, 652, long_cpuid652);
            if(active_thread[long_cpuid652])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc652_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid652/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 652 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid652]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc652_phy_pc_w))
                begin
                    if(good[long_cpuid652/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid652 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid652/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid652])
        end // if (done[652])

        if (done[653]) begin
            timeout[long_cpuid653] = 0;
            //check_bad_trap(spc653_phy_pc_w, 653, long_cpuid653);
            if(active_thread[long_cpuid653])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc653_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid653/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 653 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid653]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc653_phy_pc_w))
                begin
                    if(good[long_cpuid653/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid653 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid653/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid653])
        end // if (done[653])

        if (done[654]) begin
            timeout[long_cpuid654] = 0;
            //check_bad_trap(spc654_phy_pc_w, 654, long_cpuid654);
            if(active_thread[long_cpuid654])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc654_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid654/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 654 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid654]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc654_phy_pc_w))
                begin
                    if(good[long_cpuid654/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid654 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid654/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid654])
        end // if (done[654])

        if (done[655]) begin
            timeout[long_cpuid655] = 0;
            //check_bad_trap(spc655_phy_pc_w, 655, long_cpuid655);
            if(active_thread[long_cpuid655])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc655_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid655/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 655 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid655]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc655_phy_pc_w))
                begin
                    if(good[long_cpuid655/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid655 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid655/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid655])
        end // if (done[655])

        if (done[656]) begin
            timeout[long_cpuid656] = 0;
            //check_bad_trap(spc656_phy_pc_w, 656, long_cpuid656);
            if(active_thread[long_cpuid656])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc656_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid656/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 656 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid656]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc656_phy_pc_w))
                begin
                    if(good[long_cpuid656/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid656 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid656/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid656])
        end // if (done[656])

        if (done[657]) begin
            timeout[long_cpuid657] = 0;
            //check_bad_trap(spc657_phy_pc_w, 657, long_cpuid657);
            if(active_thread[long_cpuid657])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc657_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid657/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 657 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid657]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc657_phy_pc_w))
                begin
                    if(good[long_cpuid657/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid657 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid657/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid657])
        end // if (done[657])

        if (done[658]) begin
            timeout[long_cpuid658] = 0;
            //check_bad_trap(spc658_phy_pc_w, 658, long_cpuid658);
            if(active_thread[long_cpuid658])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc658_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid658/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 658 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid658]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc658_phy_pc_w))
                begin
                    if(good[long_cpuid658/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid658 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid658/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid658])
        end // if (done[658])

        if (done[659]) begin
            timeout[long_cpuid659] = 0;
            //check_bad_trap(spc659_phy_pc_w, 659, long_cpuid659);
            if(active_thread[long_cpuid659])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc659_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid659/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 659 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid659]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc659_phy_pc_w))
                begin
                    if(good[long_cpuid659/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid659 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid659/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid659])
        end // if (done[659])

        if (done[660]) begin
            timeout[long_cpuid660] = 0;
            //check_bad_trap(spc660_phy_pc_w, 660, long_cpuid660);
            if(active_thread[long_cpuid660])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc660_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid660/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 660 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid660]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc660_phy_pc_w))
                begin
                    if(good[long_cpuid660/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid660 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid660/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid660])
        end // if (done[660])

        if (done[661]) begin
            timeout[long_cpuid661] = 0;
            //check_bad_trap(spc661_phy_pc_w, 661, long_cpuid661);
            if(active_thread[long_cpuid661])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc661_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid661/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 661 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid661]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc661_phy_pc_w))
                begin
                    if(good[long_cpuid661/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid661 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid661/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid661])
        end // if (done[661])

        if (done[662]) begin
            timeout[long_cpuid662] = 0;
            //check_bad_trap(spc662_phy_pc_w, 662, long_cpuid662);
            if(active_thread[long_cpuid662])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc662_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid662/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 662 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid662]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc662_phy_pc_w))
                begin
                    if(good[long_cpuid662/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid662 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid662/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid662])
        end // if (done[662])

        if (done[663]) begin
            timeout[long_cpuid663] = 0;
            //check_bad_trap(spc663_phy_pc_w, 663, long_cpuid663);
            if(active_thread[long_cpuid663])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc663_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid663/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 663 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid663]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc663_phy_pc_w))
                begin
                    if(good[long_cpuid663/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid663 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid663/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid663])
        end // if (done[663])

        if (done[664]) begin
            timeout[long_cpuid664] = 0;
            //check_bad_trap(spc664_phy_pc_w, 664, long_cpuid664);
            if(active_thread[long_cpuid664])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc664_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid664/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 664 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid664]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc664_phy_pc_w))
                begin
                    if(good[long_cpuid664/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid664 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid664/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid664])
        end // if (done[664])

        if (done[665]) begin
            timeout[long_cpuid665] = 0;
            //check_bad_trap(spc665_phy_pc_w, 665, long_cpuid665);
            if(active_thread[long_cpuid665])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc665_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid665/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 665 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid665]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc665_phy_pc_w))
                begin
                    if(good[long_cpuid665/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid665 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid665/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid665])
        end // if (done[665])

        if (done[666]) begin
            timeout[long_cpuid666] = 0;
            //check_bad_trap(spc666_phy_pc_w, 666, long_cpuid666);
            if(active_thread[long_cpuid666])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc666_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid666/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 666 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid666]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc666_phy_pc_w))
                begin
                    if(good[long_cpuid666/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid666 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid666/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid666])
        end // if (done[666])

        if (done[667]) begin
            timeout[long_cpuid667] = 0;
            //check_bad_trap(spc667_phy_pc_w, 667, long_cpuid667);
            if(active_thread[long_cpuid667])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc667_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid667/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 667 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid667]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc667_phy_pc_w))
                begin
                    if(good[long_cpuid667/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid667 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid667/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid667])
        end // if (done[667])

        if (done[668]) begin
            timeout[long_cpuid668] = 0;
            //check_bad_trap(spc668_phy_pc_w, 668, long_cpuid668);
            if(active_thread[long_cpuid668])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc668_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid668/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 668 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid668]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc668_phy_pc_w))
                begin
                    if(good[long_cpuid668/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid668 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid668/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid668])
        end // if (done[668])

        if (done[669]) begin
            timeout[long_cpuid669] = 0;
            //check_bad_trap(spc669_phy_pc_w, 669, long_cpuid669);
            if(active_thread[long_cpuid669])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc669_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid669/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 669 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid669]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc669_phy_pc_w))
                begin
                    if(good[long_cpuid669/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid669 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid669/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid669])
        end // if (done[669])

        if (done[670]) begin
            timeout[long_cpuid670] = 0;
            //check_bad_trap(spc670_phy_pc_w, 670, long_cpuid670);
            if(active_thread[long_cpuid670])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc670_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid670/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 670 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid670]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc670_phy_pc_w))
                begin
                    if(good[long_cpuid670/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid670 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid670/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid670])
        end // if (done[670])

        if (done[671]) begin
            timeout[long_cpuid671] = 0;
            //check_bad_trap(spc671_phy_pc_w, 671, long_cpuid671);
            if(active_thread[long_cpuid671])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc671_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid671/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 671 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid671]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc671_phy_pc_w))
                begin
                    if(good[long_cpuid671/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid671 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid671/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid671])
        end // if (done[671])

        if (done[672]) begin
            timeout[long_cpuid672] = 0;
            //check_bad_trap(spc672_phy_pc_w, 672, long_cpuid672);
            if(active_thread[long_cpuid672])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc672_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid672/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 672 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid672]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc672_phy_pc_w))
                begin
                    if(good[long_cpuid672/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid672 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid672/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid672])
        end // if (done[672])

        if (done[673]) begin
            timeout[long_cpuid673] = 0;
            //check_bad_trap(spc673_phy_pc_w, 673, long_cpuid673);
            if(active_thread[long_cpuid673])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc673_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid673/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 673 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid673]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc673_phy_pc_w))
                begin
                    if(good[long_cpuid673/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid673 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid673/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid673])
        end // if (done[673])

        if (done[674]) begin
            timeout[long_cpuid674] = 0;
            //check_bad_trap(spc674_phy_pc_w, 674, long_cpuid674);
            if(active_thread[long_cpuid674])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc674_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid674/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 674 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid674]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc674_phy_pc_w))
                begin
                    if(good[long_cpuid674/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid674 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid674/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid674])
        end // if (done[674])

        if (done[675]) begin
            timeout[long_cpuid675] = 0;
            //check_bad_trap(spc675_phy_pc_w, 675, long_cpuid675);
            if(active_thread[long_cpuid675])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc675_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid675/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 675 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid675]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc675_phy_pc_w))
                begin
                    if(good[long_cpuid675/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid675 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid675/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid675])
        end // if (done[675])

        if (done[676]) begin
            timeout[long_cpuid676] = 0;
            //check_bad_trap(spc676_phy_pc_w, 676, long_cpuid676);
            if(active_thread[long_cpuid676])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc676_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid676/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 676 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid676]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc676_phy_pc_w))
                begin
                    if(good[long_cpuid676/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid676 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid676/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid676])
        end // if (done[676])

        if (done[677]) begin
            timeout[long_cpuid677] = 0;
            //check_bad_trap(spc677_phy_pc_w, 677, long_cpuid677);
            if(active_thread[long_cpuid677])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc677_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid677/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 677 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid677]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc677_phy_pc_w))
                begin
                    if(good[long_cpuid677/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid677 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid677/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid677])
        end // if (done[677])

        if (done[678]) begin
            timeout[long_cpuid678] = 0;
            //check_bad_trap(spc678_phy_pc_w, 678, long_cpuid678);
            if(active_thread[long_cpuid678])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc678_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid678/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 678 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid678]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc678_phy_pc_w))
                begin
                    if(good[long_cpuid678/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid678 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid678/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid678])
        end // if (done[678])

        if (done[679]) begin
            timeout[long_cpuid679] = 0;
            //check_bad_trap(spc679_phy_pc_w, 679, long_cpuid679);
            if(active_thread[long_cpuid679])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc679_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid679/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 679 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid679]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc679_phy_pc_w))
                begin
                    if(good[long_cpuid679/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid679 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid679/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid679])
        end // if (done[679])

        if (done[680]) begin
            timeout[long_cpuid680] = 0;
            //check_bad_trap(spc680_phy_pc_w, 680, long_cpuid680);
            if(active_thread[long_cpuid680])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc680_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid680/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 680 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid680]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc680_phy_pc_w))
                begin
                    if(good[long_cpuid680/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid680 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid680/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid680])
        end // if (done[680])

        if (done[681]) begin
            timeout[long_cpuid681] = 0;
            //check_bad_trap(spc681_phy_pc_w, 681, long_cpuid681);
            if(active_thread[long_cpuid681])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc681_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid681/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 681 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid681]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc681_phy_pc_w))
                begin
                    if(good[long_cpuid681/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid681 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid681/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid681])
        end // if (done[681])

        if (done[682]) begin
            timeout[long_cpuid682] = 0;
            //check_bad_trap(spc682_phy_pc_w, 682, long_cpuid682);
            if(active_thread[long_cpuid682])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc682_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid682/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 682 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid682]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc682_phy_pc_w))
                begin
                    if(good[long_cpuid682/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid682 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid682/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid682])
        end // if (done[682])

        if (done[683]) begin
            timeout[long_cpuid683] = 0;
            //check_bad_trap(spc683_phy_pc_w, 683, long_cpuid683);
            if(active_thread[long_cpuid683])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc683_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid683/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 683 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid683]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc683_phy_pc_w))
                begin
                    if(good[long_cpuid683/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid683 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid683/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid683])
        end // if (done[683])

        if (done[684]) begin
            timeout[long_cpuid684] = 0;
            //check_bad_trap(spc684_phy_pc_w, 684, long_cpuid684);
            if(active_thread[long_cpuid684])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc684_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid684/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 684 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid684]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc684_phy_pc_w))
                begin
                    if(good[long_cpuid684/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid684 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid684/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid684])
        end // if (done[684])

        if (done[685]) begin
            timeout[long_cpuid685] = 0;
            //check_bad_trap(spc685_phy_pc_w, 685, long_cpuid685);
            if(active_thread[long_cpuid685])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc685_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid685/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 685 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid685]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc685_phy_pc_w))
                begin
                    if(good[long_cpuid685/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid685 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid685/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid685])
        end // if (done[685])

        if (done[686]) begin
            timeout[long_cpuid686] = 0;
            //check_bad_trap(spc686_phy_pc_w, 686, long_cpuid686);
            if(active_thread[long_cpuid686])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc686_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid686/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 686 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid686]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc686_phy_pc_w))
                begin
                    if(good[long_cpuid686/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid686 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid686/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid686])
        end // if (done[686])

        if (done[687]) begin
            timeout[long_cpuid687] = 0;
            //check_bad_trap(spc687_phy_pc_w, 687, long_cpuid687);
            if(active_thread[long_cpuid687])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc687_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid687/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 687 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid687]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc687_phy_pc_w))
                begin
                    if(good[long_cpuid687/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid687 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid687/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid687])
        end // if (done[687])

        if (done[688]) begin
            timeout[long_cpuid688] = 0;
            //check_bad_trap(spc688_phy_pc_w, 688, long_cpuid688);
            if(active_thread[long_cpuid688])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc688_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid688/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 688 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid688]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc688_phy_pc_w))
                begin
                    if(good[long_cpuid688/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid688 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid688/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid688])
        end // if (done[688])

        if (done[689]) begin
            timeout[long_cpuid689] = 0;
            //check_bad_trap(spc689_phy_pc_w, 689, long_cpuid689);
            if(active_thread[long_cpuid689])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc689_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid689/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 689 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid689]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc689_phy_pc_w))
                begin
                    if(good[long_cpuid689/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid689 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid689/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid689])
        end // if (done[689])

        if (done[690]) begin
            timeout[long_cpuid690] = 0;
            //check_bad_trap(spc690_phy_pc_w, 690, long_cpuid690);
            if(active_thread[long_cpuid690])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc690_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid690/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 690 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid690]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc690_phy_pc_w))
                begin
                    if(good[long_cpuid690/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid690 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid690/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid690])
        end // if (done[690])

        if (done[691]) begin
            timeout[long_cpuid691] = 0;
            //check_bad_trap(spc691_phy_pc_w, 691, long_cpuid691);
            if(active_thread[long_cpuid691])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc691_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid691/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 691 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid691]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc691_phy_pc_w))
                begin
                    if(good[long_cpuid691/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid691 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid691/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid691])
        end // if (done[691])

        if (done[692]) begin
            timeout[long_cpuid692] = 0;
            //check_bad_trap(spc692_phy_pc_w, 692, long_cpuid692);
            if(active_thread[long_cpuid692])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc692_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid692/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 692 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid692]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc692_phy_pc_w))
                begin
                    if(good[long_cpuid692/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid692 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid692/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid692])
        end // if (done[692])

        if (done[693]) begin
            timeout[long_cpuid693] = 0;
            //check_bad_trap(spc693_phy_pc_w, 693, long_cpuid693);
            if(active_thread[long_cpuid693])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc693_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid693/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 693 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid693]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc693_phy_pc_w))
                begin
                    if(good[long_cpuid693/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid693 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid693/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid693])
        end // if (done[693])

        if (done[694]) begin
            timeout[long_cpuid694] = 0;
            //check_bad_trap(spc694_phy_pc_w, 694, long_cpuid694);
            if(active_thread[long_cpuid694])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc694_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid694/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 694 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid694]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc694_phy_pc_w))
                begin
                    if(good[long_cpuid694/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid694 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid694/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid694])
        end // if (done[694])

        if (done[695]) begin
            timeout[long_cpuid695] = 0;
            //check_bad_trap(spc695_phy_pc_w, 695, long_cpuid695);
            if(active_thread[long_cpuid695])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc695_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid695/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 695 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid695]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc695_phy_pc_w))
                begin
                    if(good[long_cpuid695/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid695 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid695/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid695])
        end // if (done[695])

        if (done[696]) begin
            timeout[long_cpuid696] = 0;
            //check_bad_trap(spc696_phy_pc_w, 696, long_cpuid696);
            if(active_thread[long_cpuid696])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc696_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid696/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 696 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid696]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc696_phy_pc_w))
                begin
                    if(good[long_cpuid696/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid696 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid696/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid696])
        end // if (done[696])

        if (done[697]) begin
            timeout[long_cpuid697] = 0;
            //check_bad_trap(spc697_phy_pc_w, 697, long_cpuid697);
            if(active_thread[long_cpuid697])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc697_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid697/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 697 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid697]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc697_phy_pc_w))
                begin
                    if(good[long_cpuid697/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid697 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid697/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid697])
        end // if (done[697])

        if (done[698]) begin
            timeout[long_cpuid698] = 0;
            //check_bad_trap(spc698_phy_pc_w, 698, long_cpuid698);
            if(active_thread[long_cpuid698])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc698_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid698/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 698 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid698]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc698_phy_pc_w))
                begin
                    if(good[long_cpuid698/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid698 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid698/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid698])
        end // if (done[698])

        if (done[699]) begin
            timeout[long_cpuid699] = 0;
            //check_bad_trap(spc699_phy_pc_w, 699, long_cpuid699);
            if(active_thread[long_cpuid699])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc699_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid699/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 699 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid699]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc699_phy_pc_w))
                begin
                    if(good[long_cpuid699/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid699 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid699/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid699])
        end // if (done[699])

        if (done[700]) begin
            timeout[long_cpuid700] = 0;
            //check_bad_trap(spc700_phy_pc_w, 700, long_cpuid700);
            if(active_thread[long_cpuid700])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc700_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid700/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 700 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid700]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc700_phy_pc_w))
                begin
                    if(good[long_cpuid700/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid700 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid700/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid700])
        end // if (done[700])

        if (done[701]) begin
            timeout[long_cpuid701] = 0;
            //check_bad_trap(spc701_phy_pc_w, 701, long_cpuid701);
            if(active_thread[long_cpuid701])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc701_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid701/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 701 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid701]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc701_phy_pc_w))
                begin
                    if(good[long_cpuid701/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid701 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid701/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid701])
        end // if (done[701])

        if (done[702]) begin
            timeout[long_cpuid702] = 0;
            //check_bad_trap(spc702_phy_pc_w, 702, long_cpuid702);
            if(active_thread[long_cpuid702])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc702_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid702/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 702 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid702]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc702_phy_pc_w))
                begin
                    if(good[long_cpuid702/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid702 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid702/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid702])
        end // if (done[702])

        if (done[703]) begin
            timeout[long_cpuid703] = 0;
            //check_bad_trap(spc703_phy_pc_w, 703, long_cpuid703);
            if(active_thread[long_cpuid703])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc703_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid703/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 703 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid703]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc703_phy_pc_w))
                begin
                    if(good[long_cpuid703/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid703 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid703/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid703])
        end // if (done[703])

        if (done[704]) begin
            timeout[long_cpuid704] = 0;
            //check_bad_trap(spc704_phy_pc_w, 704, long_cpuid704);
            if(active_thread[long_cpuid704])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc704_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid704/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 704 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid704]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc704_phy_pc_w))
                begin
                    if(good[long_cpuid704/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid704 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid704/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid704])
        end // if (done[704])

        if (done[705]) begin
            timeout[long_cpuid705] = 0;
            //check_bad_trap(spc705_phy_pc_w, 705, long_cpuid705);
            if(active_thread[long_cpuid705])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc705_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid705/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 705 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid705]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc705_phy_pc_w))
                begin
                    if(good[long_cpuid705/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid705 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid705/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid705])
        end // if (done[705])

        if (done[706]) begin
            timeout[long_cpuid706] = 0;
            //check_bad_trap(spc706_phy_pc_w, 706, long_cpuid706);
            if(active_thread[long_cpuid706])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc706_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid706/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 706 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid706]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc706_phy_pc_w))
                begin
                    if(good[long_cpuid706/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid706 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid706/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid706])
        end // if (done[706])

        if (done[707]) begin
            timeout[long_cpuid707] = 0;
            //check_bad_trap(spc707_phy_pc_w, 707, long_cpuid707);
            if(active_thread[long_cpuid707])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc707_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid707/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 707 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid707]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc707_phy_pc_w))
                begin
                    if(good[long_cpuid707/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid707 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid707/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid707])
        end // if (done[707])

        if (done[708]) begin
            timeout[long_cpuid708] = 0;
            //check_bad_trap(spc708_phy_pc_w, 708, long_cpuid708);
            if(active_thread[long_cpuid708])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc708_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid708/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 708 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid708]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc708_phy_pc_w))
                begin
                    if(good[long_cpuid708/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid708 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid708/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid708])
        end // if (done[708])

        if (done[709]) begin
            timeout[long_cpuid709] = 0;
            //check_bad_trap(spc709_phy_pc_w, 709, long_cpuid709);
            if(active_thread[long_cpuid709])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc709_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid709/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 709 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid709]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc709_phy_pc_w))
                begin
                    if(good[long_cpuid709/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid709 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid709/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid709])
        end // if (done[709])

        if (done[710]) begin
            timeout[long_cpuid710] = 0;
            //check_bad_trap(spc710_phy_pc_w, 710, long_cpuid710);
            if(active_thread[long_cpuid710])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc710_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid710/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 710 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid710]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc710_phy_pc_w))
                begin
                    if(good[long_cpuid710/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid710 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid710/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid710])
        end // if (done[710])

        if (done[711]) begin
            timeout[long_cpuid711] = 0;
            //check_bad_trap(spc711_phy_pc_w, 711, long_cpuid711);
            if(active_thread[long_cpuid711])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc711_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid711/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 711 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid711]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc711_phy_pc_w))
                begin
                    if(good[long_cpuid711/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid711 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid711/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid711])
        end // if (done[711])

        if (done[712]) begin
            timeout[long_cpuid712] = 0;
            //check_bad_trap(spc712_phy_pc_w, 712, long_cpuid712);
            if(active_thread[long_cpuid712])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc712_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid712/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 712 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid712]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc712_phy_pc_w))
                begin
                    if(good[long_cpuid712/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid712 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid712/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid712])
        end // if (done[712])

        if (done[713]) begin
            timeout[long_cpuid713] = 0;
            //check_bad_trap(spc713_phy_pc_w, 713, long_cpuid713);
            if(active_thread[long_cpuid713])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc713_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid713/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 713 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid713]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc713_phy_pc_w))
                begin
                    if(good[long_cpuid713/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid713 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid713/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid713])
        end // if (done[713])

        if (done[714]) begin
            timeout[long_cpuid714] = 0;
            //check_bad_trap(spc714_phy_pc_w, 714, long_cpuid714);
            if(active_thread[long_cpuid714])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc714_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid714/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 714 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid714]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc714_phy_pc_w))
                begin
                    if(good[long_cpuid714/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid714 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid714/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid714])
        end // if (done[714])

        if (done[715]) begin
            timeout[long_cpuid715] = 0;
            //check_bad_trap(spc715_phy_pc_w, 715, long_cpuid715);
            if(active_thread[long_cpuid715])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc715_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid715/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 715 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid715]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc715_phy_pc_w))
                begin
                    if(good[long_cpuid715/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid715 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid715/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid715])
        end // if (done[715])

        if (done[716]) begin
            timeout[long_cpuid716] = 0;
            //check_bad_trap(spc716_phy_pc_w, 716, long_cpuid716);
            if(active_thread[long_cpuid716])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc716_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid716/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 716 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid716]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc716_phy_pc_w))
                begin
                    if(good[long_cpuid716/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid716 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid716/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid716])
        end // if (done[716])

        if (done[717]) begin
            timeout[long_cpuid717] = 0;
            //check_bad_trap(spc717_phy_pc_w, 717, long_cpuid717);
            if(active_thread[long_cpuid717])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc717_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid717/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 717 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid717]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc717_phy_pc_w))
                begin
                    if(good[long_cpuid717/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid717 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid717/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid717])
        end // if (done[717])

        if (done[718]) begin
            timeout[long_cpuid718] = 0;
            //check_bad_trap(spc718_phy_pc_w, 718, long_cpuid718);
            if(active_thread[long_cpuid718])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc718_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid718/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 718 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid718]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc718_phy_pc_w))
                begin
                    if(good[long_cpuid718/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid718 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid718/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid718])
        end // if (done[718])

        if (done[719]) begin
            timeout[long_cpuid719] = 0;
            //check_bad_trap(spc719_phy_pc_w, 719, long_cpuid719);
            if(active_thread[long_cpuid719])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc719_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid719/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 719 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid719]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc719_phy_pc_w))
                begin
                    if(good[long_cpuid719/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid719 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid719/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid719])
        end // if (done[719])

        if (done[720]) begin
            timeout[long_cpuid720] = 0;
            //check_bad_trap(spc720_phy_pc_w, 720, long_cpuid720);
            if(active_thread[long_cpuid720])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc720_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid720/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 720 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid720]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc720_phy_pc_w))
                begin
                    if(good[long_cpuid720/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid720 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid720/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid720])
        end // if (done[720])

        if (done[721]) begin
            timeout[long_cpuid721] = 0;
            //check_bad_trap(spc721_phy_pc_w, 721, long_cpuid721);
            if(active_thread[long_cpuid721])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc721_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid721/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 721 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid721]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc721_phy_pc_w))
                begin
                    if(good[long_cpuid721/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid721 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid721/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid721])
        end // if (done[721])

        if (done[722]) begin
            timeout[long_cpuid722] = 0;
            //check_bad_trap(spc722_phy_pc_w, 722, long_cpuid722);
            if(active_thread[long_cpuid722])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc722_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid722/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 722 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid722]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc722_phy_pc_w))
                begin
                    if(good[long_cpuid722/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid722 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid722/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid722])
        end // if (done[722])

        if (done[723]) begin
            timeout[long_cpuid723] = 0;
            //check_bad_trap(spc723_phy_pc_w, 723, long_cpuid723);
            if(active_thread[long_cpuid723])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc723_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid723/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 723 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid723]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc723_phy_pc_w))
                begin
                    if(good[long_cpuid723/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid723 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid723/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid723])
        end // if (done[723])

        if (done[724]) begin
            timeout[long_cpuid724] = 0;
            //check_bad_trap(spc724_phy_pc_w, 724, long_cpuid724);
            if(active_thread[long_cpuid724])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc724_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid724/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 724 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid724]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc724_phy_pc_w))
                begin
                    if(good[long_cpuid724/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid724 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid724/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid724])
        end // if (done[724])

        if (done[725]) begin
            timeout[long_cpuid725] = 0;
            //check_bad_trap(spc725_phy_pc_w, 725, long_cpuid725);
            if(active_thread[long_cpuid725])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc725_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid725/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 725 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid725]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc725_phy_pc_w))
                begin
                    if(good[long_cpuid725/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid725 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid725/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid725])
        end // if (done[725])

        if (done[726]) begin
            timeout[long_cpuid726] = 0;
            //check_bad_trap(spc726_phy_pc_w, 726, long_cpuid726);
            if(active_thread[long_cpuid726])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc726_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid726/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 726 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid726]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc726_phy_pc_w))
                begin
                    if(good[long_cpuid726/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid726 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid726/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid726])
        end // if (done[726])

        if (done[727]) begin
            timeout[long_cpuid727] = 0;
            //check_bad_trap(spc727_phy_pc_w, 727, long_cpuid727);
            if(active_thread[long_cpuid727])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc727_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid727/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 727 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid727]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc727_phy_pc_w))
                begin
                    if(good[long_cpuid727/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid727 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid727/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid727])
        end // if (done[727])

        if (done[728]) begin
            timeout[long_cpuid728] = 0;
            //check_bad_trap(spc728_phy_pc_w, 728, long_cpuid728);
            if(active_thread[long_cpuid728])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc728_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid728/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 728 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid728]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc728_phy_pc_w))
                begin
                    if(good[long_cpuid728/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid728 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid728/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid728])
        end // if (done[728])

        if (done[729]) begin
            timeout[long_cpuid729] = 0;
            //check_bad_trap(spc729_phy_pc_w, 729, long_cpuid729);
            if(active_thread[long_cpuid729])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc729_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid729/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 729 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid729]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc729_phy_pc_w))
                begin
                    if(good[long_cpuid729/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid729 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid729/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid729])
        end // if (done[729])

        if (done[730]) begin
            timeout[long_cpuid730] = 0;
            //check_bad_trap(spc730_phy_pc_w, 730, long_cpuid730);
            if(active_thread[long_cpuid730])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc730_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid730/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 730 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid730]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc730_phy_pc_w))
                begin
                    if(good[long_cpuid730/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid730 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid730/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid730])
        end // if (done[730])

        if (done[731]) begin
            timeout[long_cpuid731] = 0;
            //check_bad_trap(spc731_phy_pc_w, 731, long_cpuid731);
            if(active_thread[long_cpuid731])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc731_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid731/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 731 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid731]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc731_phy_pc_w))
                begin
                    if(good[long_cpuid731/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid731 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid731/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid731])
        end // if (done[731])

        if (done[732]) begin
            timeout[long_cpuid732] = 0;
            //check_bad_trap(spc732_phy_pc_w, 732, long_cpuid732);
            if(active_thread[long_cpuid732])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc732_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid732/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 732 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid732]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc732_phy_pc_w))
                begin
                    if(good[long_cpuid732/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid732 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid732/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid732])
        end // if (done[732])

        if (done[733]) begin
            timeout[long_cpuid733] = 0;
            //check_bad_trap(spc733_phy_pc_w, 733, long_cpuid733);
            if(active_thread[long_cpuid733])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc733_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid733/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 733 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid733]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc733_phy_pc_w))
                begin
                    if(good[long_cpuid733/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid733 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid733/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid733])
        end // if (done[733])

        if (done[734]) begin
            timeout[long_cpuid734] = 0;
            //check_bad_trap(spc734_phy_pc_w, 734, long_cpuid734);
            if(active_thread[long_cpuid734])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc734_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid734/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 734 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid734]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc734_phy_pc_w))
                begin
                    if(good[long_cpuid734/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid734 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid734/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid734])
        end // if (done[734])

        if (done[735]) begin
            timeout[long_cpuid735] = 0;
            //check_bad_trap(spc735_phy_pc_w, 735, long_cpuid735);
            if(active_thread[long_cpuid735])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc735_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid735/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 735 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid735]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc735_phy_pc_w))
                begin
                    if(good[long_cpuid735/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid735 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid735/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid735])
        end // if (done[735])

        if (done[736]) begin
            timeout[long_cpuid736] = 0;
            //check_bad_trap(spc736_phy_pc_w, 736, long_cpuid736);
            if(active_thread[long_cpuid736])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc736_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid736/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 736 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid736]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc736_phy_pc_w))
                begin
                    if(good[long_cpuid736/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid736 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid736/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid736])
        end // if (done[736])

        if (done[737]) begin
            timeout[long_cpuid737] = 0;
            //check_bad_trap(spc737_phy_pc_w, 737, long_cpuid737);
            if(active_thread[long_cpuid737])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc737_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid737/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 737 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid737]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc737_phy_pc_w))
                begin
                    if(good[long_cpuid737/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid737 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid737/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid737])
        end // if (done[737])

        if (done[738]) begin
            timeout[long_cpuid738] = 0;
            //check_bad_trap(spc738_phy_pc_w, 738, long_cpuid738);
            if(active_thread[long_cpuid738])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc738_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid738/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 738 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid738]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc738_phy_pc_w))
                begin
                    if(good[long_cpuid738/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid738 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid738/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid738])
        end // if (done[738])

        if (done[739]) begin
            timeout[long_cpuid739] = 0;
            //check_bad_trap(spc739_phy_pc_w, 739, long_cpuid739);
            if(active_thread[long_cpuid739])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc739_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid739/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 739 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid739]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc739_phy_pc_w))
                begin
                    if(good[long_cpuid739/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid739 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid739/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid739])
        end // if (done[739])

        if (done[740]) begin
            timeout[long_cpuid740] = 0;
            //check_bad_trap(spc740_phy_pc_w, 740, long_cpuid740);
            if(active_thread[long_cpuid740])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc740_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid740/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 740 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid740]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc740_phy_pc_w))
                begin
                    if(good[long_cpuid740/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid740 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid740/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid740])
        end // if (done[740])

        if (done[741]) begin
            timeout[long_cpuid741] = 0;
            //check_bad_trap(spc741_phy_pc_w, 741, long_cpuid741);
            if(active_thread[long_cpuid741])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc741_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid741/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 741 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid741]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc741_phy_pc_w))
                begin
                    if(good[long_cpuid741/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid741 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid741/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid741])
        end // if (done[741])

        if (done[742]) begin
            timeout[long_cpuid742] = 0;
            //check_bad_trap(spc742_phy_pc_w, 742, long_cpuid742);
            if(active_thread[long_cpuid742])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc742_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid742/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 742 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid742]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc742_phy_pc_w))
                begin
                    if(good[long_cpuid742/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid742 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid742/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid742])
        end // if (done[742])

        if (done[743]) begin
            timeout[long_cpuid743] = 0;
            //check_bad_trap(spc743_phy_pc_w, 743, long_cpuid743);
            if(active_thread[long_cpuid743])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc743_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid743/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 743 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid743]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc743_phy_pc_w))
                begin
                    if(good[long_cpuid743/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid743 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid743/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid743])
        end // if (done[743])

        if (done[744]) begin
            timeout[long_cpuid744] = 0;
            //check_bad_trap(spc744_phy_pc_w, 744, long_cpuid744);
            if(active_thread[long_cpuid744])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc744_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid744/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 744 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid744]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc744_phy_pc_w))
                begin
                    if(good[long_cpuid744/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid744 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid744/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid744])
        end // if (done[744])

        if (done[745]) begin
            timeout[long_cpuid745] = 0;
            //check_bad_trap(spc745_phy_pc_w, 745, long_cpuid745);
            if(active_thread[long_cpuid745])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc745_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid745/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 745 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid745]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc745_phy_pc_w))
                begin
                    if(good[long_cpuid745/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid745 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid745/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid745])
        end // if (done[745])

        if (done[746]) begin
            timeout[long_cpuid746] = 0;
            //check_bad_trap(spc746_phy_pc_w, 746, long_cpuid746);
            if(active_thread[long_cpuid746])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc746_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid746/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 746 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid746]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc746_phy_pc_w))
                begin
                    if(good[long_cpuid746/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid746 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid746/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid746])
        end // if (done[746])

        if (done[747]) begin
            timeout[long_cpuid747] = 0;
            //check_bad_trap(spc747_phy_pc_w, 747, long_cpuid747);
            if(active_thread[long_cpuid747])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc747_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid747/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 747 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid747]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc747_phy_pc_w))
                begin
                    if(good[long_cpuid747/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid747 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid747/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid747])
        end // if (done[747])

        if (done[748]) begin
            timeout[long_cpuid748] = 0;
            //check_bad_trap(spc748_phy_pc_w, 748, long_cpuid748);
            if(active_thread[long_cpuid748])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc748_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid748/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 748 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid748]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc748_phy_pc_w))
                begin
                    if(good[long_cpuid748/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid748 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid748/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid748])
        end // if (done[748])

        if (done[749]) begin
            timeout[long_cpuid749] = 0;
            //check_bad_trap(spc749_phy_pc_w, 749, long_cpuid749);
            if(active_thread[long_cpuid749])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc749_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid749/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 749 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid749]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc749_phy_pc_w))
                begin
                    if(good[long_cpuid749/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid749 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid749/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid749])
        end // if (done[749])

        if (done[750]) begin
            timeout[long_cpuid750] = 0;
            //check_bad_trap(spc750_phy_pc_w, 750, long_cpuid750);
            if(active_thread[long_cpuid750])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc750_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid750/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 750 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid750]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc750_phy_pc_w))
                begin
                    if(good[long_cpuid750/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid750 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid750/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid750])
        end // if (done[750])

        if (done[751]) begin
            timeout[long_cpuid751] = 0;
            //check_bad_trap(spc751_phy_pc_w, 751, long_cpuid751);
            if(active_thread[long_cpuid751])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc751_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid751/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 751 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid751]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc751_phy_pc_w))
                begin
                    if(good[long_cpuid751/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid751 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid751/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid751])
        end // if (done[751])

        if (done[752]) begin
            timeout[long_cpuid752] = 0;
            //check_bad_trap(spc752_phy_pc_w, 752, long_cpuid752);
            if(active_thread[long_cpuid752])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc752_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid752/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 752 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid752]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc752_phy_pc_w))
                begin
                    if(good[long_cpuid752/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid752 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid752/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid752])
        end // if (done[752])

        if (done[753]) begin
            timeout[long_cpuid753] = 0;
            //check_bad_trap(spc753_phy_pc_w, 753, long_cpuid753);
            if(active_thread[long_cpuid753])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc753_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid753/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 753 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid753]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc753_phy_pc_w))
                begin
                    if(good[long_cpuid753/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid753 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid753/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid753])
        end // if (done[753])

        if (done[754]) begin
            timeout[long_cpuid754] = 0;
            //check_bad_trap(spc754_phy_pc_w, 754, long_cpuid754);
            if(active_thread[long_cpuid754])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc754_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid754/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 754 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid754]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc754_phy_pc_w))
                begin
                    if(good[long_cpuid754/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid754 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid754/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid754])
        end // if (done[754])

        if (done[755]) begin
            timeout[long_cpuid755] = 0;
            //check_bad_trap(spc755_phy_pc_w, 755, long_cpuid755);
            if(active_thread[long_cpuid755])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc755_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid755/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 755 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid755]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc755_phy_pc_w))
                begin
                    if(good[long_cpuid755/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid755 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid755/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid755])
        end // if (done[755])

        if (done[756]) begin
            timeout[long_cpuid756] = 0;
            //check_bad_trap(spc756_phy_pc_w, 756, long_cpuid756);
            if(active_thread[long_cpuid756])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc756_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid756/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 756 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid756]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc756_phy_pc_w))
                begin
                    if(good[long_cpuid756/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid756 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid756/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid756])
        end // if (done[756])

        if (done[757]) begin
            timeout[long_cpuid757] = 0;
            //check_bad_trap(spc757_phy_pc_w, 757, long_cpuid757);
            if(active_thread[long_cpuid757])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc757_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid757/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 757 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid757]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc757_phy_pc_w))
                begin
                    if(good[long_cpuid757/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid757 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid757/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid757])
        end // if (done[757])

        if (done[758]) begin
            timeout[long_cpuid758] = 0;
            //check_bad_trap(spc758_phy_pc_w, 758, long_cpuid758);
            if(active_thread[long_cpuid758])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc758_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid758/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 758 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid758]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc758_phy_pc_w))
                begin
                    if(good[long_cpuid758/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid758 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid758/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid758])
        end // if (done[758])

        if (done[759]) begin
            timeout[long_cpuid759] = 0;
            //check_bad_trap(spc759_phy_pc_w, 759, long_cpuid759);
            if(active_thread[long_cpuid759])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc759_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid759/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 759 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid759]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc759_phy_pc_w))
                begin
                    if(good[long_cpuid759/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid759 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid759/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid759])
        end // if (done[759])

        if (done[760]) begin
            timeout[long_cpuid760] = 0;
            //check_bad_trap(spc760_phy_pc_w, 760, long_cpuid760);
            if(active_thread[long_cpuid760])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc760_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid760/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 760 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid760]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc760_phy_pc_w))
                begin
                    if(good[long_cpuid760/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid760 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid760/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid760])
        end // if (done[760])

        if (done[761]) begin
            timeout[long_cpuid761] = 0;
            //check_bad_trap(spc761_phy_pc_w, 761, long_cpuid761);
            if(active_thread[long_cpuid761])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc761_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid761/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 761 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid761]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc761_phy_pc_w))
                begin
                    if(good[long_cpuid761/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid761 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid761/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid761])
        end // if (done[761])

        if (done[762]) begin
            timeout[long_cpuid762] = 0;
            //check_bad_trap(spc762_phy_pc_w, 762, long_cpuid762);
            if(active_thread[long_cpuid762])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc762_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid762/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 762 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid762]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc762_phy_pc_w))
                begin
                    if(good[long_cpuid762/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid762 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid762/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid762])
        end // if (done[762])

        if (done[763]) begin
            timeout[long_cpuid763] = 0;
            //check_bad_trap(spc763_phy_pc_w, 763, long_cpuid763);
            if(active_thread[long_cpuid763])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc763_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid763/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 763 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid763]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc763_phy_pc_w))
                begin
                    if(good[long_cpuid763/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid763 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid763/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid763])
        end // if (done[763])

        if (done[764]) begin
            timeout[long_cpuid764] = 0;
            //check_bad_trap(spc764_phy_pc_w, 764, long_cpuid764);
            if(active_thread[long_cpuid764])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc764_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid764/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 764 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid764]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc764_phy_pc_w))
                begin
                    if(good[long_cpuid764/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid764 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid764/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid764])
        end // if (done[764])

        if (done[765]) begin
            timeout[long_cpuid765] = 0;
            //check_bad_trap(spc765_phy_pc_w, 765, long_cpuid765);
            if(active_thread[long_cpuid765])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc765_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid765/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 765 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid765]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc765_phy_pc_w))
                begin
                    if(good[long_cpuid765/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid765 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid765/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid765])
        end // if (done[765])

        if (done[766]) begin
            timeout[long_cpuid766] = 0;
            //check_bad_trap(spc766_phy_pc_w, 766, long_cpuid766);
            if(active_thread[long_cpuid766])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc766_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid766/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 766 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid766]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc766_phy_pc_w))
                begin
                    if(good[long_cpuid766/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid766 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid766/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid766])
        end // if (done[766])

        if (done[767]) begin
            timeout[long_cpuid767] = 0;
            //check_bad_trap(spc767_phy_pc_w, 767, long_cpuid767);
            if(active_thread[long_cpuid767])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc767_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid767/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 767 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid767]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc767_phy_pc_w))
                begin
                    if(good[long_cpuid767/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid767 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid767/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid767])
        end // if (done[767])

        if (done[768]) begin
            timeout[long_cpuid768] = 0;
            //check_bad_trap(spc768_phy_pc_w, 768, long_cpuid768);
            if(active_thread[long_cpuid768])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc768_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid768/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 768 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid768]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc768_phy_pc_w))
                begin
                    if(good[long_cpuid768/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid768 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid768/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid768])
        end // if (done[768])

        if (done[769]) begin
            timeout[long_cpuid769] = 0;
            //check_bad_trap(spc769_phy_pc_w, 769, long_cpuid769);
            if(active_thread[long_cpuid769])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc769_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid769/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 769 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid769]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc769_phy_pc_w))
                begin
                    if(good[long_cpuid769/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid769 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid769/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid769])
        end // if (done[769])

        if (done[770]) begin
            timeout[long_cpuid770] = 0;
            //check_bad_trap(spc770_phy_pc_w, 770, long_cpuid770);
            if(active_thread[long_cpuid770])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc770_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid770/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 770 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid770]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc770_phy_pc_w))
                begin
                    if(good[long_cpuid770/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid770 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid770/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid770])
        end // if (done[770])

        if (done[771]) begin
            timeout[long_cpuid771] = 0;
            //check_bad_trap(spc771_phy_pc_w, 771, long_cpuid771);
            if(active_thread[long_cpuid771])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc771_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid771/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 771 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid771]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc771_phy_pc_w))
                begin
                    if(good[long_cpuid771/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid771 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid771/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid771])
        end // if (done[771])

        if (done[772]) begin
            timeout[long_cpuid772] = 0;
            //check_bad_trap(spc772_phy_pc_w, 772, long_cpuid772);
            if(active_thread[long_cpuid772])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc772_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid772/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 772 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid772]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc772_phy_pc_w))
                begin
                    if(good[long_cpuid772/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid772 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid772/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid772])
        end // if (done[772])

        if (done[773]) begin
            timeout[long_cpuid773] = 0;
            //check_bad_trap(spc773_phy_pc_w, 773, long_cpuid773);
            if(active_thread[long_cpuid773])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc773_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid773/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 773 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid773]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc773_phy_pc_w))
                begin
                    if(good[long_cpuid773/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid773 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid773/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid773])
        end // if (done[773])

        if (done[774]) begin
            timeout[long_cpuid774] = 0;
            //check_bad_trap(spc774_phy_pc_w, 774, long_cpuid774);
            if(active_thread[long_cpuid774])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc774_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid774/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 774 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid774]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc774_phy_pc_w))
                begin
                    if(good[long_cpuid774/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid774 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid774/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid774])
        end // if (done[774])

        if (done[775]) begin
            timeout[long_cpuid775] = 0;
            //check_bad_trap(spc775_phy_pc_w, 775, long_cpuid775);
            if(active_thread[long_cpuid775])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc775_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid775/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 775 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid775]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc775_phy_pc_w))
                begin
                    if(good[long_cpuid775/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid775 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid775/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid775])
        end // if (done[775])

        if (done[776]) begin
            timeout[long_cpuid776] = 0;
            //check_bad_trap(spc776_phy_pc_w, 776, long_cpuid776);
            if(active_thread[long_cpuid776])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc776_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid776/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 776 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid776]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc776_phy_pc_w))
                begin
                    if(good[long_cpuid776/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid776 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid776/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid776])
        end // if (done[776])

        if (done[777]) begin
            timeout[long_cpuid777] = 0;
            //check_bad_trap(spc777_phy_pc_w, 777, long_cpuid777);
            if(active_thread[long_cpuid777])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc777_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid777/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 777 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid777]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc777_phy_pc_w))
                begin
                    if(good[long_cpuid777/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid777 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid777/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid777])
        end // if (done[777])

        if (done[778]) begin
            timeout[long_cpuid778] = 0;
            //check_bad_trap(spc778_phy_pc_w, 778, long_cpuid778);
            if(active_thread[long_cpuid778])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc778_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid778/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 778 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid778]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc778_phy_pc_w))
                begin
                    if(good[long_cpuid778/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid778 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid778/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid778])
        end // if (done[778])

        if (done[779]) begin
            timeout[long_cpuid779] = 0;
            //check_bad_trap(spc779_phy_pc_w, 779, long_cpuid779);
            if(active_thread[long_cpuid779])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc779_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid779/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 779 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid779]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc779_phy_pc_w))
                begin
                    if(good[long_cpuid779/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid779 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid779/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid779])
        end // if (done[779])

        if (done[780]) begin
            timeout[long_cpuid780] = 0;
            //check_bad_trap(spc780_phy_pc_w, 780, long_cpuid780);
            if(active_thread[long_cpuid780])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc780_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid780/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 780 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid780]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc780_phy_pc_w))
                begin
                    if(good[long_cpuid780/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid780 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid780/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid780])
        end // if (done[780])

        if (done[781]) begin
            timeout[long_cpuid781] = 0;
            //check_bad_trap(spc781_phy_pc_w, 781, long_cpuid781);
            if(active_thread[long_cpuid781])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc781_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid781/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 781 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid781]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc781_phy_pc_w))
                begin
                    if(good[long_cpuid781/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid781 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid781/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid781])
        end // if (done[781])

        if (done[782]) begin
            timeout[long_cpuid782] = 0;
            //check_bad_trap(spc782_phy_pc_w, 782, long_cpuid782);
            if(active_thread[long_cpuid782])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc782_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid782/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 782 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid782]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc782_phy_pc_w))
                begin
                    if(good[long_cpuid782/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid782 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid782/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid782])
        end // if (done[782])

        if (done[783]) begin
            timeout[long_cpuid783] = 0;
            //check_bad_trap(spc783_phy_pc_w, 783, long_cpuid783);
            if(active_thread[long_cpuid783])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc783_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid783/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 783 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid783]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc783_phy_pc_w))
                begin
                    if(good[long_cpuid783/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid783 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid783/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid783])
        end // if (done[783])

        if (done[784]) begin
            timeout[long_cpuid784] = 0;
            //check_bad_trap(spc784_phy_pc_w, 784, long_cpuid784);
            if(active_thread[long_cpuid784])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc784_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid784/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 784 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid784]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc784_phy_pc_w))
                begin
                    if(good[long_cpuid784/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid784 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid784/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid784])
        end // if (done[784])

        if (done[785]) begin
            timeout[long_cpuid785] = 0;
            //check_bad_trap(spc785_phy_pc_w, 785, long_cpuid785);
            if(active_thread[long_cpuid785])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc785_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid785/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 785 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid785]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc785_phy_pc_w))
                begin
                    if(good[long_cpuid785/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid785 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid785/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid785])
        end // if (done[785])

        if (done[786]) begin
            timeout[long_cpuid786] = 0;
            //check_bad_trap(spc786_phy_pc_w, 786, long_cpuid786);
            if(active_thread[long_cpuid786])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc786_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid786/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 786 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid786]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc786_phy_pc_w))
                begin
                    if(good[long_cpuid786/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid786 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid786/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid786])
        end // if (done[786])

        if (done[787]) begin
            timeout[long_cpuid787] = 0;
            //check_bad_trap(spc787_phy_pc_w, 787, long_cpuid787);
            if(active_thread[long_cpuid787])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc787_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid787/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 787 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid787]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc787_phy_pc_w))
                begin
                    if(good[long_cpuid787/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid787 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid787/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid787])
        end // if (done[787])

        if (done[788]) begin
            timeout[long_cpuid788] = 0;
            //check_bad_trap(spc788_phy_pc_w, 788, long_cpuid788);
            if(active_thread[long_cpuid788])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc788_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid788/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 788 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid788]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc788_phy_pc_w))
                begin
                    if(good[long_cpuid788/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid788 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid788/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid788])
        end // if (done[788])

        if (done[789]) begin
            timeout[long_cpuid789] = 0;
            //check_bad_trap(spc789_phy_pc_w, 789, long_cpuid789);
            if(active_thread[long_cpuid789])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc789_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid789/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 789 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid789]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc789_phy_pc_w))
                begin
                    if(good[long_cpuid789/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid789 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid789/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid789])
        end // if (done[789])

        if (done[790]) begin
            timeout[long_cpuid790] = 0;
            //check_bad_trap(spc790_phy_pc_w, 790, long_cpuid790);
            if(active_thread[long_cpuid790])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc790_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid790/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 790 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid790]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc790_phy_pc_w))
                begin
                    if(good[long_cpuid790/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid790 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid790/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid790])
        end // if (done[790])

        if (done[791]) begin
            timeout[long_cpuid791] = 0;
            //check_bad_trap(spc791_phy_pc_w, 791, long_cpuid791);
            if(active_thread[long_cpuid791])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc791_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid791/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 791 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid791]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc791_phy_pc_w))
                begin
                    if(good[long_cpuid791/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid791 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid791/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid791])
        end // if (done[791])

        if (done[792]) begin
            timeout[long_cpuid792] = 0;
            //check_bad_trap(spc792_phy_pc_w, 792, long_cpuid792);
            if(active_thread[long_cpuid792])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc792_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid792/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 792 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid792]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc792_phy_pc_w))
                begin
                    if(good[long_cpuid792/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid792 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid792/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid792])
        end // if (done[792])

        if (done[793]) begin
            timeout[long_cpuid793] = 0;
            //check_bad_trap(spc793_phy_pc_w, 793, long_cpuid793);
            if(active_thread[long_cpuid793])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc793_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid793/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 793 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid793]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc793_phy_pc_w))
                begin
                    if(good[long_cpuid793/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid793 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid793/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid793])
        end // if (done[793])

        if (done[794]) begin
            timeout[long_cpuid794] = 0;
            //check_bad_trap(spc794_phy_pc_w, 794, long_cpuid794);
            if(active_thread[long_cpuid794])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc794_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid794/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 794 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid794]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc794_phy_pc_w))
                begin
                    if(good[long_cpuid794/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid794 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid794/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid794])
        end // if (done[794])

        if (done[795]) begin
            timeout[long_cpuid795] = 0;
            //check_bad_trap(spc795_phy_pc_w, 795, long_cpuid795);
            if(active_thread[long_cpuid795])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc795_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid795/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 795 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid795]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc795_phy_pc_w))
                begin
                    if(good[long_cpuid795/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid795 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid795/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid795])
        end // if (done[795])

        if (done[796]) begin
            timeout[long_cpuid796] = 0;
            //check_bad_trap(spc796_phy_pc_w, 796, long_cpuid796);
            if(active_thread[long_cpuid796])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc796_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid796/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 796 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid796]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc796_phy_pc_w))
                begin
                    if(good[long_cpuid796/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid796 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid796/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid796])
        end // if (done[796])

        if (done[797]) begin
            timeout[long_cpuid797] = 0;
            //check_bad_trap(spc797_phy_pc_w, 797, long_cpuid797);
            if(active_thread[long_cpuid797])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc797_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid797/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 797 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid797]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc797_phy_pc_w))
                begin
                    if(good[long_cpuid797/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid797 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid797/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid797])
        end // if (done[797])

        if (done[798]) begin
            timeout[long_cpuid798] = 0;
            //check_bad_trap(spc798_phy_pc_w, 798, long_cpuid798);
            if(active_thread[long_cpuid798])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc798_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid798/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 798 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid798]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc798_phy_pc_w))
                begin
                    if(good[long_cpuid798/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid798 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid798/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid798])
        end // if (done[798])

        if (done[799]) begin
            timeout[long_cpuid799] = 0;
            //check_bad_trap(spc799_phy_pc_w, 799, long_cpuid799);
            if(active_thread[long_cpuid799])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc799_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid799/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 799 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid799]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc799_phy_pc_w))
                begin
                    if(good[long_cpuid799/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid799 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid799/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid799])
        end // if (done[799])

        if (done[800]) begin
            timeout[long_cpuid800] = 0;
            //check_bad_trap(spc800_phy_pc_w, 800, long_cpuid800);
            if(active_thread[long_cpuid800])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc800_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid800/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 800 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid800]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc800_phy_pc_w))
                begin
                    if(good[long_cpuid800/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid800 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid800/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid800])
        end // if (done[800])

        if (done[801]) begin
            timeout[long_cpuid801] = 0;
            //check_bad_trap(spc801_phy_pc_w, 801, long_cpuid801);
            if(active_thread[long_cpuid801])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc801_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid801/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 801 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid801]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc801_phy_pc_w))
                begin
                    if(good[long_cpuid801/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid801 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid801/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid801])
        end // if (done[801])

        if (done[802]) begin
            timeout[long_cpuid802] = 0;
            //check_bad_trap(spc802_phy_pc_w, 802, long_cpuid802);
            if(active_thread[long_cpuid802])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc802_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid802/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 802 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid802]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc802_phy_pc_w))
                begin
                    if(good[long_cpuid802/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid802 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid802/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid802])
        end // if (done[802])

        if (done[803]) begin
            timeout[long_cpuid803] = 0;
            //check_bad_trap(spc803_phy_pc_w, 803, long_cpuid803);
            if(active_thread[long_cpuid803])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc803_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid803/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 803 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid803]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc803_phy_pc_w))
                begin
                    if(good[long_cpuid803/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid803 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid803/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid803])
        end // if (done[803])

        if (done[804]) begin
            timeout[long_cpuid804] = 0;
            //check_bad_trap(spc804_phy_pc_w, 804, long_cpuid804);
            if(active_thread[long_cpuid804])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc804_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid804/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 804 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid804]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc804_phy_pc_w))
                begin
                    if(good[long_cpuid804/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid804 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid804/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid804])
        end // if (done[804])

        if (done[805]) begin
            timeout[long_cpuid805] = 0;
            //check_bad_trap(spc805_phy_pc_w, 805, long_cpuid805);
            if(active_thread[long_cpuid805])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc805_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid805/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 805 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid805]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc805_phy_pc_w))
                begin
                    if(good[long_cpuid805/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid805 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid805/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid805])
        end // if (done[805])

        if (done[806]) begin
            timeout[long_cpuid806] = 0;
            //check_bad_trap(spc806_phy_pc_w, 806, long_cpuid806);
            if(active_thread[long_cpuid806])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc806_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid806/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 806 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid806]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc806_phy_pc_w))
                begin
                    if(good[long_cpuid806/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid806 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid806/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid806])
        end // if (done[806])

        if (done[807]) begin
            timeout[long_cpuid807] = 0;
            //check_bad_trap(spc807_phy_pc_w, 807, long_cpuid807);
            if(active_thread[long_cpuid807])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc807_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid807/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 807 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid807]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc807_phy_pc_w))
                begin
                    if(good[long_cpuid807/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid807 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid807/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid807])
        end // if (done[807])

        if (done[808]) begin
            timeout[long_cpuid808] = 0;
            //check_bad_trap(spc808_phy_pc_w, 808, long_cpuid808);
            if(active_thread[long_cpuid808])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc808_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid808/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 808 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid808]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc808_phy_pc_w))
                begin
                    if(good[long_cpuid808/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid808 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid808/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid808])
        end // if (done[808])

        if (done[809]) begin
            timeout[long_cpuid809] = 0;
            //check_bad_trap(spc809_phy_pc_w, 809, long_cpuid809);
            if(active_thread[long_cpuid809])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc809_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid809/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 809 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid809]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc809_phy_pc_w))
                begin
                    if(good[long_cpuid809/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid809 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid809/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid809])
        end // if (done[809])

        if (done[810]) begin
            timeout[long_cpuid810] = 0;
            //check_bad_trap(spc810_phy_pc_w, 810, long_cpuid810);
            if(active_thread[long_cpuid810])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc810_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid810/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 810 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid810]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc810_phy_pc_w))
                begin
                    if(good[long_cpuid810/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid810 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid810/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid810])
        end // if (done[810])

        if (done[811]) begin
            timeout[long_cpuid811] = 0;
            //check_bad_trap(spc811_phy_pc_w, 811, long_cpuid811);
            if(active_thread[long_cpuid811])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc811_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid811/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 811 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid811]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc811_phy_pc_w))
                begin
                    if(good[long_cpuid811/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid811 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid811/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid811])
        end // if (done[811])

        if (done[812]) begin
            timeout[long_cpuid812] = 0;
            //check_bad_trap(spc812_phy_pc_w, 812, long_cpuid812);
            if(active_thread[long_cpuid812])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc812_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid812/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 812 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid812]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc812_phy_pc_w))
                begin
                    if(good[long_cpuid812/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid812 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid812/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid812])
        end // if (done[812])

        if (done[813]) begin
            timeout[long_cpuid813] = 0;
            //check_bad_trap(spc813_phy_pc_w, 813, long_cpuid813);
            if(active_thread[long_cpuid813])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc813_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid813/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 813 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid813]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc813_phy_pc_w))
                begin
                    if(good[long_cpuid813/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid813 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid813/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid813])
        end // if (done[813])

        if (done[814]) begin
            timeout[long_cpuid814] = 0;
            //check_bad_trap(spc814_phy_pc_w, 814, long_cpuid814);
            if(active_thread[long_cpuid814])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc814_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid814/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 814 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid814]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc814_phy_pc_w))
                begin
                    if(good[long_cpuid814/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid814 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid814/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid814])
        end // if (done[814])

        if (done[815]) begin
            timeout[long_cpuid815] = 0;
            //check_bad_trap(spc815_phy_pc_w, 815, long_cpuid815);
            if(active_thread[long_cpuid815])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc815_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid815/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 815 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid815]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc815_phy_pc_w))
                begin
                    if(good[long_cpuid815/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid815 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid815/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid815])
        end // if (done[815])

        if (done[816]) begin
            timeout[long_cpuid816] = 0;
            //check_bad_trap(spc816_phy_pc_w, 816, long_cpuid816);
            if(active_thread[long_cpuid816])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc816_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid816/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 816 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid816]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc816_phy_pc_w))
                begin
                    if(good[long_cpuid816/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid816 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid816/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid816])
        end // if (done[816])

        if (done[817]) begin
            timeout[long_cpuid817] = 0;
            //check_bad_trap(spc817_phy_pc_w, 817, long_cpuid817);
            if(active_thread[long_cpuid817])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc817_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid817/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 817 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid817]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc817_phy_pc_w))
                begin
                    if(good[long_cpuid817/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid817 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid817/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid817])
        end // if (done[817])

        if (done[818]) begin
            timeout[long_cpuid818] = 0;
            //check_bad_trap(spc818_phy_pc_w, 818, long_cpuid818);
            if(active_thread[long_cpuid818])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc818_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid818/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 818 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid818]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc818_phy_pc_w))
                begin
                    if(good[long_cpuid818/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid818 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid818/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid818])
        end // if (done[818])

        if (done[819]) begin
            timeout[long_cpuid819] = 0;
            //check_bad_trap(spc819_phy_pc_w, 819, long_cpuid819);
            if(active_thread[long_cpuid819])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc819_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid819/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 819 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid819]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc819_phy_pc_w))
                begin
                    if(good[long_cpuid819/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid819 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid819/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid819])
        end // if (done[819])

        if (done[820]) begin
            timeout[long_cpuid820] = 0;
            //check_bad_trap(spc820_phy_pc_w, 820, long_cpuid820);
            if(active_thread[long_cpuid820])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc820_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid820/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 820 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid820]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc820_phy_pc_w))
                begin
                    if(good[long_cpuid820/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid820 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid820/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid820])
        end // if (done[820])

        if (done[821]) begin
            timeout[long_cpuid821] = 0;
            //check_bad_trap(spc821_phy_pc_w, 821, long_cpuid821);
            if(active_thread[long_cpuid821])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc821_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid821/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 821 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid821]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc821_phy_pc_w))
                begin
                    if(good[long_cpuid821/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid821 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid821/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid821])
        end // if (done[821])

        if (done[822]) begin
            timeout[long_cpuid822] = 0;
            //check_bad_trap(spc822_phy_pc_w, 822, long_cpuid822);
            if(active_thread[long_cpuid822])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc822_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid822/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 822 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid822]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc822_phy_pc_w))
                begin
                    if(good[long_cpuid822/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid822 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid822/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid822])
        end // if (done[822])

        if (done[823]) begin
            timeout[long_cpuid823] = 0;
            //check_bad_trap(spc823_phy_pc_w, 823, long_cpuid823);
            if(active_thread[long_cpuid823])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc823_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid823/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 823 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid823]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc823_phy_pc_w))
                begin
                    if(good[long_cpuid823/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid823 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid823/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid823])
        end // if (done[823])

        if (done[824]) begin
            timeout[long_cpuid824] = 0;
            //check_bad_trap(spc824_phy_pc_w, 824, long_cpuid824);
            if(active_thread[long_cpuid824])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc824_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid824/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 824 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid824]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc824_phy_pc_w))
                begin
                    if(good[long_cpuid824/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid824 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid824/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid824])
        end // if (done[824])

        if (done[825]) begin
            timeout[long_cpuid825] = 0;
            //check_bad_trap(spc825_phy_pc_w, 825, long_cpuid825);
            if(active_thread[long_cpuid825])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc825_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid825/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 825 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid825]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc825_phy_pc_w))
                begin
                    if(good[long_cpuid825/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid825 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid825/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid825])
        end // if (done[825])

        if (done[826]) begin
            timeout[long_cpuid826] = 0;
            //check_bad_trap(spc826_phy_pc_w, 826, long_cpuid826);
            if(active_thread[long_cpuid826])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc826_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid826/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 826 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid826]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc826_phy_pc_w))
                begin
                    if(good[long_cpuid826/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid826 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid826/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid826])
        end // if (done[826])

        if (done[827]) begin
            timeout[long_cpuid827] = 0;
            //check_bad_trap(spc827_phy_pc_w, 827, long_cpuid827);
            if(active_thread[long_cpuid827])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc827_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid827/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 827 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid827]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc827_phy_pc_w))
                begin
                    if(good[long_cpuid827/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid827 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid827/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid827])
        end // if (done[827])

        if (done[828]) begin
            timeout[long_cpuid828] = 0;
            //check_bad_trap(spc828_phy_pc_w, 828, long_cpuid828);
            if(active_thread[long_cpuid828])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc828_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid828/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 828 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid828]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc828_phy_pc_w))
                begin
                    if(good[long_cpuid828/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid828 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid828/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid828])
        end // if (done[828])

        if (done[829]) begin
            timeout[long_cpuid829] = 0;
            //check_bad_trap(spc829_phy_pc_w, 829, long_cpuid829);
            if(active_thread[long_cpuid829])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc829_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid829/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 829 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid829]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc829_phy_pc_w))
                begin
                    if(good[long_cpuid829/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid829 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid829/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid829])
        end // if (done[829])

        if (done[830]) begin
            timeout[long_cpuid830] = 0;
            //check_bad_trap(spc830_phy_pc_w, 830, long_cpuid830);
            if(active_thread[long_cpuid830])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc830_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid830/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 830 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid830]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc830_phy_pc_w))
                begin
                    if(good[long_cpuid830/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid830 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid830/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid830])
        end // if (done[830])

        if (done[831]) begin
            timeout[long_cpuid831] = 0;
            //check_bad_trap(spc831_phy_pc_w, 831, long_cpuid831);
            if(active_thread[long_cpuid831])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc831_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid831/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 831 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid831]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc831_phy_pc_w))
                begin
                    if(good[long_cpuid831/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid831 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid831/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid831])
        end // if (done[831])

        if (done[832]) begin
            timeout[long_cpuid832] = 0;
            //check_bad_trap(spc832_phy_pc_w, 832, long_cpuid832);
            if(active_thread[long_cpuid832])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc832_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid832/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 832 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid832]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc832_phy_pc_w))
                begin
                    if(good[long_cpuid832/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid832 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid832/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid832])
        end // if (done[832])

        if (done[833]) begin
            timeout[long_cpuid833] = 0;
            //check_bad_trap(spc833_phy_pc_w, 833, long_cpuid833);
            if(active_thread[long_cpuid833])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc833_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid833/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 833 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid833]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc833_phy_pc_w))
                begin
                    if(good[long_cpuid833/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid833 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid833/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid833])
        end // if (done[833])

        if (done[834]) begin
            timeout[long_cpuid834] = 0;
            //check_bad_trap(spc834_phy_pc_w, 834, long_cpuid834);
            if(active_thread[long_cpuid834])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc834_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid834/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 834 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid834]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc834_phy_pc_w))
                begin
                    if(good[long_cpuid834/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid834 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid834/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid834])
        end // if (done[834])

        if (done[835]) begin
            timeout[long_cpuid835] = 0;
            //check_bad_trap(spc835_phy_pc_w, 835, long_cpuid835);
            if(active_thread[long_cpuid835])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc835_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid835/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 835 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid835]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc835_phy_pc_w))
                begin
                    if(good[long_cpuid835/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid835 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid835/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid835])
        end // if (done[835])

        if (done[836]) begin
            timeout[long_cpuid836] = 0;
            //check_bad_trap(spc836_phy_pc_w, 836, long_cpuid836);
            if(active_thread[long_cpuid836])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc836_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid836/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 836 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid836]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc836_phy_pc_w))
                begin
                    if(good[long_cpuid836/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid836 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid836/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid836])
        end // if (done[836])

        if (done[837]) begin
            timeout[long_cpuid837] = 0;
            //check_bad_trap(spc837_phy_pc_w, 837, long_cpuid837);
            if(active_thread[long_cpuid837])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc837_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid837/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 837 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid837]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc837_phy_pc_w))
                begin
                    if(good[long_cpuid837/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid837 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid837/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid837])
        end // if (done[837])

        if (done[838]) begin
            timeout[long_cpuid838] = 0;
            //check_bad_trap(spc838_phy_pc_w, 838, long_cpuid838);
            if(active_thread[long_cpuid838])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc838_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid838/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 838 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid838]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc838_phy_pc_w))
                begin
                    if(good[long_cpuid838/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid838 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid838/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid838])
        end // if (done[838])

        if (done[839]) begin
            timeout[long_cpuid839] = 0;
            //check_bad_trap(spc839_phy_pc_w, 839, long_cpuid839);
            if(active_thread[long_cpuid839])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc839_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid839/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 839 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid839]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc839_phy_pc_w))
                begin
                    if(good[long_cpuid839/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid839 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid839/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid839])
        end // if (done[839])

        if (done[840]) begin
            timeout[long_cpuid840] = 0;
            //check_bad_trap(spc840_phy_pc_w, 840, long_cpuid840);
            if(active_thread[long_cpuid840])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc840_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid840/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 840 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid840]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc840_phy_pc_w))
                begin
                    if(good[long_cpuid840/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid840 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid840/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid840])
        end // if (done[840])

        if (done[841]) begin
            timeout[long_cpuid841] = 0;
            //check_bad_trap(spc841_phy_pc_w, 841, long_cpuid841);
            if(active_thread[long_cpuid841])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc841_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid841/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 841 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid841]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc841_phy_pc_w))
                begin
                    if(good[long_cpuid841/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid841 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid841/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid841])
        end // if (done[841])

        if (done[842]) begin
            timeout[long_cpuid842] = 0;
            //check_bad_trap(spc842_phy_pc_w, 842, long_cpuid842);
            if(active_thread[long_cpuid842])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc842_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid842/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 842 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid842]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc842_phy_pc_w))
                begin
                    if(good[long_cpuid842/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid842 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid842/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid842])
        end // if (done[842])

        if (done[843]) begin
            timeout[long_cpuid843] = 0;
            //check_bad_trap(spc843_phy_pc_w, 843, long_cpuid843);
            if(active_thread[long_cpuid843])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc843_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid843/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 843 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid843]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc843_phy_pc_w))
                begin
                    if(good[long_cpuid843/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid843 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid843/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid843])
        end // if (done[843])

        if (done[844]) begin
            timeout[long_cpuid844] = 0;
            //check_bad_trap(spc844_phy_pc_w, 844, long_cpuid844);
            if(active_thread[long_cpuid844])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc844_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid844/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 844 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid844]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc844_phy_pc_w))
                begin
                    if(good[long_cpuid844/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid844 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid844/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid844])
        end // if (done[844])

        if (done[845]) begin
            timeout[long_cpuid845] = 0;
            //check_bad_trap(spc845_phy_pc_w, 845, long_cpuid845);
            if(active_thread[long_cpuid845])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc845_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid845/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 845 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid845]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc845_phy_pc_w))
                begin
                    if(good[long_cpuid845/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid845 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid845/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid845])
        end // if (done[845])

        if (done[846]) begin
            timeout[long_cpuid846] = 0;
            //check_bad_trap(spc846_phy_pc_w, 846, long_cpuid846);
            if(active_thread[long_cpuid846])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc846_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid846/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 846 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid846]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc846_phy_pc_w))
                begin
                    if(good[long_cpuid846/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid846 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid846/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid846])
        end // if (done[846])

        if (done[847]) begin
            timeout[long_cpuid847] = 0;
            //check_bad_trap(spc847_phy_pc_w, 847, long_cpuid847);
            if(active_thread[long_cpuid847])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc847_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid847/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 847 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid847]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc847_phy_pc_w))
                begin
                    if(good[long_cpuid847/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid847 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid847/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid847])
        end // if (done[847])

        if (done[848]) begin
            timeout[long_cpuid848] = 0;
            //check_bad_trap(spc848_phy_pc_w, 848, long_cpuid848);
            if(active_thread[long_cpuid848])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc848_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid848/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 848 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid848]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc848_phy_pc_w))
                begin
                    if(good[long_cpuid848/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid848 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid848/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid848])
        end // if (done[848])

        if (done[849]) begin
            timeout[long_cpuid849] = 0;
            //check_bad_trap(spc849_phy_pc_w, 849, long_cpuid849);
            if(active_thread[long_cpuid849])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc849_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid849/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 849 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid849]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc849_phy_pc_w))
                begin
                    if(good[long_cpuid849/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid849 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid849/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid849])
        end // if (done[849])

        if (done[850]) begin
            timeout[long_cpuid850] = 0;
            //check_bad_trap(spc850_phy_pc_w, 850, long_cpuid850);
            if(active_thread[long_cpuid850])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc850_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid850/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 850 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid850]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc850_phy_pc_w))
                begin
                    if(good[long_cpuid850/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid850 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid850/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid850])
        end // if (done[850])

        if (done[851]) begin
            timeout[long_cpuid851] = 0;
            //check_bad_trap(spc851_phy_pc_w, 851, long_cpuid851);
            if(active_thread[long_cpuid851])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc851_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid851/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 851 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid851]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc851_phy_pc_w))
                begin
                    if(good[long_cpuid851/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid851 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid851/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid851])
        end // if (done[851])

        if (done[852]) begin
            timeout[long_cpuid852] = 0;
            //check_bad_trap(spc852_phy_pc_w, 852, long_cpuid852);
            if(active_thread[long_cpuid852])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc852_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid852/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 852 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid852]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc852_phy_pc_w))
                begin
                    if(good[long_cpuid852/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid852 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid852/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid852])
        end // if (done[852])

        if (done[853]) begin
            timeout[long_cpuid853] = 0;
            //check_bad_trap(spc853_phy_pc_w, 853, long_cpuid853);
            if(active_thread[long_cpuid853])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc853_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid853/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 853 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid853]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc853_phy_pc_w))
                begin
                    if(good[long_cpuid853/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid853 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid853/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid853])
        end // if (done[853])

        if (done[854]) begin
            timeout[long_cpuid854] = 0;
            //check_bad_trap(spc854_phy_pc_w, 854, long_cpuid854);
            if(active_thread[long_cpuid854])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc854_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid854/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 854 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid854]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc854_phy_pc_w))
                begin
                    if(good[long_cpuid854/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid854 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid854/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid854])
        end // if (done[854])

        if (done[855]) begin
            timeout[long_cpuid855] = 0;
            //check_bad_trap(spc855_phy_pc_w, 855, long_cpuid855);
            if(active_thread[long_cpuid855])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc855_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid855/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 855 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid855]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc855_phy_pc_w))
                begin
                    if(good[long_cpuid855/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid855 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid855/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid855])
        end // if (done[855])

        if (done[856]) begin
            timeout[long_cpuid856] = 0;
            //check_bad_trap(spc856_phy_pc_w, 856, long_cpuid856);
            if(active_thread[long_cpuid856])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc856_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid856/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 856 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid856]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc856_phy_pc_w))
                begin
                    if(good[long_cpuid856/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid856 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid856/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid856])
        end // if (done[856])

        if (done[857]) begin
            timeout[long_cpuid857] = 0;
            //check_bad_trap(spc857_phy_pc_w, 857, long_cpuid857);
            if(active_thread[long_cpuid857])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc857_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid857/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 857 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid857]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc857_phy_pc_w))
                begin
                    if(good[long_cpuid857/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid857 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid857/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid857])
        end // if (done[857])

        if (done[858]) begin
            timeout[long_cpuid858] = 0;
            //check_bad_trap(spc858_phy_pc_w, 858, long_cpuid858);
            if(active_thread[long_cpuid858])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc858_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid858/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 858 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid858]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc858_phy_pc_w))
                begin
                    if(good[long_cpuid858/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid858 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid858/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid858])
        end // if (done[858])

        if (done[859]) begin
            timeout[long_cpuid859] = 0;
            //check_bad_trap(spc859_phy_pc_w, 859, long_cpuid859);
            if(active_thread[long_cpuid859])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc859_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid859/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 859 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid859]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc859_phy_pc_w))
                begin
                    if(good[long_cpuid859/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid859 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid859/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid859])
        end // if (done[859])

        if (done[860]) begin
            timeout[long_cpuid860] = 0;
            //check_bad_trap(spc860_phy_pc_w, 860, long_cpuid860);
            if(active_thread[long_cpuid860])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc860_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid860/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 860 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid860]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc860_phy_pc_w))
                begin
                    if(good[long_cpuid860/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid860 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid860/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid860])
        end // if (done[860])

        if (done[861]) begin
            timeout[long_cpuid861] = 0;
            //check_bad_trap(spc861_phy_pc_w, 861, long_cpuid861);
            if(active_thread[long_cpuid861])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc861_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid861/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 861 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid861]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc861_phy_pc_w))
                begin
                    if(good[long_cpuid861/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid861 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid861/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid861])
        end // if (done[861])

        if (done[862]) begin
            timeout[long_cpuid862] = 0;
            //check_bad_trap(spc862_phy_pc_w, 862, long_cpuid862);
            if(active_thread[long_cpuid862])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc862_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid862/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 862 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid862]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc862_phy_pc_w))
                begin
                    if(good[long_cpuid862/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid862 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid862/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid862])
        end // if (done[862])

        if (done[863]) begin
            timeout[long_cpuid863] = 0;
            //check_bad_trap(spc863_phy_pc_w, 863, long_cpuid863);
            if(active_thread[long_cpuid863])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc863_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid863/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 863 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid863]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc863_phy_pc_w))
                begin
                    if(good[long_cpuid863/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid863 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid863/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid863])
        end // if (done[863])

        if (done[864]) begin
            timeout[long_cpuid864] = 0;
            //check_bad_trap(spc864_phy_pc_w, 864, long_cpuid864);
            if(active_thread[long_cpuid864])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc864_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid864/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 864 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid864]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc864_phy_pc_w))
                begin
                    if(good[long_cpuid864/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid864 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid864/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid864])
        end // if (done[864])

        if (done[865]) begin
            timeout[long_cpuid865] = 0;
            //check_bad_trap(spc865_phy_pc_w, 865, long_cpuid865);
            if(active_thread[long_cpuid865])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc865_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid865/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 865 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid865]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc865_phy_pc_w))
                begin
                    if(good[long_cpuid865/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid865 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid865/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid865])
        end // if (done[865])

        if (done[866]) begin
            timeout[long_cpuid866] = 0;
            //check_bad_trap(spc866_phy_pc_w, 866, long_cpuid866);
            if(active_thread[long_cpuid866])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc866_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid866/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 866 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid866]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc866_phy_pc_w))
                begin
                    if(good[long_cpuid866/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid866 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid866/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid866])
        end // if (done[866])

        if (done[867]) begin
            timeout[long_cpuid867] = 0;
            //check_bad_trap(spc867_phy_pc_w, 867, long_cpuid867);
            if(active_thread[long_cpuid867])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc867_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid867/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 867 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid867]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc867_phy_pc_w))
                begin
                    if(good[long_cpuid867/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid867 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid867/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid867])
        end // if (done[867])

        if (done[868]) begin
            timeout[long_cpuid868] = 0;
            //check_bad_trap(spc868_phy_pc_w, 868, long_cpuid868);
            if(active_thread[long_cpuid868])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc868_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid868/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 868 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid868]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc868_phy_pc_w))
                begin
                    if(good[long_cpuid868/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid868 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid868/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid868])
        end // if (done[868])

        if (done[869]) begin
            timeout[long_cpuid869] = 0;
            //check_bad_trap(spc869_phy_pc_w, 869, long_cpuid869);
            if(active_thread[long_cpuid869])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc869_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid869/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 869 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid869]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc869_phy_pc_w))
                begin
                    if(good[long_cpuid869/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid869 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid869/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid869])
        end // if (done[869])

        if (done[870]) begin
            timeout[long_cpuid870] = 0;
            //check_bad_trap(spc870_phy_pc_w, 870, long_cpuid870);
            if(active_thread[long_cpuid870])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc870_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid870/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 870 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid870]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc870_phy_pc_w))
                begin
                    if(good[long_cpuid870/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid870 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid870/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid870])
        end // if (done[870])

        if (done[871]) begin
            timeout[long_cpuid871] = 0;
            //check_bad_trap(spc871_phy_pc_w, 871, long_cpuid871);
            if(active_thread[long_cpuid871])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc871_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid871/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 871 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid871]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc871_phy_pc_w))
                begin
                    if(good[long_cpuid871/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid871 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid871/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid871])
        end // if (done[871])

        if (done[872]) begin
            timeout[long_cpuid872] = 0;
            //check_bad_trap(spc872_phy_pc_w, 872, long_cpuid872);
            if(active_thread[long_cpuid872])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc872_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid872/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 872 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid872]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc872_phy_pc_w))
                begin
                    if(good[long_cpuid872/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid872 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid872/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid872])
        end // if (done[872])

        if (done[873]) begin
            timeout[long_cpuid873] = 0;
            //check_bad_trap(spc873_phy_pc_w, 873, long_cpuid873);
            if(active_thread[long_cpuid873])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc873_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid873/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 873 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid873]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc873_phy_pc_w))
                begin
                    if(good[long_cpuid873/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid873 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid873/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid873])
        end // if (done[873])

        if (done[874]) begin
            timeout[long_cpuid874] = 0;
            //check_bad_trap(spc874_phy_pc_w, 874, long_cpuid874);
            if(active_thread[long_cpuid874])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc874_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid874/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 874 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid874]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc874_phy_pc_w))
                begin
                    if(good[long_cpuid874/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid874 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid874/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid874])
        end // if (done[874])

        if (done[875]) begin
            timeout[long_cpuid875] = 0;
            //check_bad_trap(spc875_phy_pc_w, 875, long_cpuid875);
            if(active_thread[long_cpuid875])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc875_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid875/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 875 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid875]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc875_phy_pc_w))
                begin
                    if(good[long_cpuid875/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid875 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid875/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid875])
        end // if (done[875])

        if (done[876]) begin
            timeout[long_cpuid876] = 0;
            //check_bad_trap(spc876_phy_pc_w, 876, long_cpuid876);
            if(active_thread[long_cpuid876])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc876_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid876/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 876 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid876]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc876_phy_pc_w))
                begin
                    if(good[long_cpuid876/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid876 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid876/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid876])
        end // if (done[876])

        if (done[877]) begin
            timeout[long_cpuid877] = 0;
            //check_bad_trap(spc877_phy_pc_w, 877, long_cpuid877);
            if(active_thread[long_cpuid877])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc877_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid877/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 877 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid877]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc877_phy_pc_w))
                begin
                    if(good[long_cpuid877/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid877 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid877/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid877])
        end // if (done[877])

        if (done[878]) begin
            timeout[long_cpuid878] = 0;
            //check_bad_trap(spc878_phy_pc_w, 878, long_cpuid878);
            if(active_thread[long_cpuid878])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc878_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid878/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 878 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid878]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc878_phy_pc_w))
                begin
                    if(good[long_cpuid878/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid878 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid878/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid878])
        end // if (done[878])

        if (done[879]) begin
            timeout[long_cpuid879] = 0;
            //check_bad_trap(spc879_phy_pc_w, 879, long_cpuid879);
            if(active_thread[long_cpuid879])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc879_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid879/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 879 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid879]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc879_phy_pc_w))
                begin
                    if(good[long_cpuid879/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid879 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid879/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid879])
        end // if (done[879])

        if (done[880]) begin
            timeout[long_cpuid880] = 0;
            //check_bad_trap(spc880_phy_pc_w, 880, long_cpuid880);
            if(active_thread[long_cpuid880])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc880_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid880/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 880 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid880]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc880_phy_pc_w))
                begin
                    if(good[long_cpuid880/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid880 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid880/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid880])
        end // if (done[880])

        if (done[881]) begin
            timeout[long_cpuid881] = 0;
            //check_bad_trap(spc881_phy_pc_w, 881, long_cpuid881);
            if(active_thread[long_cpuid881])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc881_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid881/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 881 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid881]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc881_phy_pc_w))
                begin
                    if(good[long_cpuid881/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid881 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid881/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid881])
        end // if (done[881])

        if (done[882]) begin
            timeout[long_cpuid882] = 0;
            //check_bad_trap(spc882_phy_pc_w, 882, long_cpuid882);
            if(active_thread[long_cpuid882])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc882_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid882/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 882 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid882]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc882_phy_pc_w))
                begin
                    if(good[long_cpuid882/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid882 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid882/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid882])
        end // if (done[882])

        if (done[883]) begin
            timeout[long_cpuid883] = 0;
            //check_bad_trap(spc883_phy_pc_w, 883, long_cpuid883);
            if(active_thread[long_cpuid883])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc883_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid883/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 883 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid883]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc883_phy_pc_w))
                begin
                    if(good[long_cpuid883/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid883 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid883/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid883])
        end // if (done[883])

        if (done[884]) begin
            timeout[long_cpuid884] = 0;
            //check_bad_trap(spc884_phy_pc_w, 884, long_cpuid884);
            if(active_thread[long_cpuid884])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc884_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid884/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 884 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid884]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc884_phy_pc_w))
                begin
                    if(good[long_cpuid884/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid884 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid884/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid884])
        end // if (done[884])

        if (done[885]) begin
            timeout[long_cpuid885] = 0;
            //check_bad_trap(spc885_phy_pc_w, 885, long_cpuid885);
            if(active_thread[long_cpuid885])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc885_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid885/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 885 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid885]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc885_phy_pc_w))
                begin
                    if(good[long_cpuid885/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid885 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid885/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid885])
        end // if (done[885])

        if (done[886]) begin
            timeout[long_cpuid886] = 0;
            //check_bad_trap(spc886_phy_pc_w, 886, long_cpuid886);
            if(active_thread[long_cpuid886])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc886_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid886/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 886 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid886]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc886_phy_pc_w))
                begin
                    if(good[long_cpuid886/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid886 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid886/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid886])
        end // if (done[886])

        if (done[887]) begin
            timeout[long_cpuid887] = 0;
            //check_bad_trap(spc887_phy_pc_w, 887, long_cpuid887);
            if(active_thread[long_cpuid887])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc887_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid887/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 887 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid887]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc887_phy_pc_w))
                begin
                    if(good[long_cpuid887/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid887 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid887/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid887])
        end // if (done[887])

        if (done[888]) begin
            timeout[long_cpuid888] = 0;
            //check_bad_trap(spc888_phy_pc_w, 888, long_cpuid888);
            if(active_thread[long_cpuid888])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc888_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid888/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 888 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid888]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc888_phy_pc_w))
                begin
                    if(good[long_cpuid888/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid888 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid888/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid888])
        end // if (done[888])

        if (done[889]) begin
            timeout[long_cpuid889] = 0;
            //check_bad_trap(spc889_phy_pc_w, 889, long_cpuid889);
            if(active_thread[long_cpuid889])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc889_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid889/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 889 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid889]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc889_phy_pc_w))
                begin
                    if(good[long_cpuid889/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid889 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid889/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid889])
        end // if (done[889])

        if (done[890]) begin
            timeout[long_cpuid890] = 0;
            //check_bad_trap(spc890_phy_pc_w, 890, long_cpuid890);
            if(active_thread[long_cpuid890])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc890_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid890/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 890 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid890]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc890_phy_pc_w))
                begin
                    if(good[long_cpuid890/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid890 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid890/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid890])
        end // if (done[890])

        if (done[891]) begin
            timeout[long_cpuid891] = 0;
            //check_bad_trap(spc891_phy_pc_w, 891, long_cpuid891);
            if(active_thread[long_cpuid891])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc891_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid891/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 891 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid891]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc891_phy_pc_w))
                begin
                    if(good[long_cpuid891/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid891 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid891/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid891])
        end // if (done[891])

        if (done[892]) begin
            timeout[long_cpuid892] = 0;
            //check_bad_trap(spc892_phy_pc_w, 892, long_cpuid892);
            if(active_thread[long_cpuid892])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc892_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid892/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 892 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid892]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc892_phy_pc_w))
                begin
                    if(good[long_cpuid892/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid892 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid892/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid892])
        end // if (done[892])

        if (done[893]) begin
            timeout[long_cpuid893] = 0;
            //check_bad_trap(spc893_phy_pc_w, 893, long_cpuid893);
            if(active_thread[long_cpuid893])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc893_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid893/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 893 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid893]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc893_phy_pc_w))
                begin
                    if(good[long_cpuid893/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid893 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid893/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid893])
        end // if (done[893])

        if (done[894]) begin
            timeout[long_cpuid894] = 0;
            //check_bad_trap(spc894_phy_pc_w, 894, long_cpuid894);
            if(active_thread[long_cpuid894])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc894_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid894/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 894 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid894]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc894_phy_pc_w))
                begin
                    if(good[long_cpuid894/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid894 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid894/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid894])
        end // if (done[894])

        if (done[895]) begin
            timeout[long_cpuid895] = 0;
            //check_bad_trap(spc895_phy_pc_w, 895, long_cpuid895);
            if(active_thread[long_cpuid895])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc895_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid895/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 895 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid895]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc895_phy_pc_w))
                begin
                    if(good[long_cpuid895/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid895 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid895/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid895])
        end // if (done[895])

        if (done[896]) begin
            timeout[long_cpuid896] = 0;
            //check_bad_trap(spc896_phy_pc_w, 896, long_cpuid896);
            if(active_thread[long_cpuid896])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc896_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid896/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 896 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid896]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc896_phy_pc_w))
                begin
                    if(good[long_cpuid896/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid896 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid896/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid896])
        end // if (done[896])

        if (done[897]) begin
            timeout[long_cpuid897] = 0;
            //check_bad_trap(spc897_phy_pc_w, 897, long_cpuid897);
            if(active_thread[long_cpuid897])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc897_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid897/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 897 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid897]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc897_phy_pc_w))
                begin
                    if(good[long_cpuid897/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid897 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid897/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid897])
        end // if (done[897])

        if (done[898]) begin
            timeout[long_cpuid898] = 0;
            //check_bad_trap(spc898_phy_pc_w, 898, long_cpuid898);
            if(active_thread[long_cpuid898])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc898_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid898/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 898 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid898]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc898_phy_pc_w))
                begin
                    if(good[long_cpuid898/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid898 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid898/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid898])
        end // if (done[898])

        if (done[899]) begin
            timeout[long_cpuid899] = 0;
            //check_bad_trap(spc899_phy_pc_w, 899, long_cpuid899);
            if(active_thread[long_cpuid899])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc899_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid899/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 899 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid899]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc899_phy_pc_w))
                begin
                    if(good[long_cpuid899/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid899 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid899/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid899])
        end // if (done[899])

        if (done[900]) begin
            timeout[long_cpuid900] = 0;
            //check_bad_trap(spc900_phy_pc_w, 900, long_cpuid900);
            if(active_thread[long_cpuid900])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc900_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid900/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 900 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid900]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc900_phy_pc_w))
                begin
                    if(good[long_cpuid900/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid900 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid900/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid900])
        end // if (done[900])

        if (done[901]) begin
            timeout[long_cpuid901] = 0;
            //check_bad_trap(spc901_phy_pc_w, 901, long_cpuid901);
            if(active_thread[long_cpuid901])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc901_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid901/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 901 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid901]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc901_phy_pc_w))
                begin
                    if(good[long_cpuid901/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid901 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid901/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid901])
        end // if (done[901])

        if (done[902]) begin
            timeout[long_cpuid902] = 0;
            //check_bad_trap(spc902_phy_pc_w, 902, long_cpuid902);
            if(active_thread[long_cpuid902])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc902_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid902/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 902 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid902]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc902_phy_pc_w))
                begin
                    if(good[long_cpuid902/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid902 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid902/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid902])
        end // if (done[902])

        if (done[903]) begin
            timeout[long_cpuid903] = 0;
            //check_bad_trap(spc903_phy_pc_w, 903, long_cpuid903);
            if(active_thread[long_cpuid903])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc903_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid903/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 903 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid903]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc903_phy_pc_w))
                begin
                    if(good[long_cpuid903/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid903 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid903/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid903])
        end // if (done[903])

        if (done[904]) begin
            timeout[long_cpuid904] = 0;
            //check_bad_trap(spc904_phy_pc_w, 904, long_cpuid904);
            if(active_thread[long_cpuid904])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc904_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid904/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 904 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid904]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc904_phy_pc_w))
                begin
                    if(good[long_cpuid904/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid904 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid904/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid904])
        end // if (done[904])

        if (done[905]) begin
            timeout[long_cpuid905] = 0;
            //check_bad_trap(spc905_phy_pc_w, 905, long_cpuid905);
            if(active_thread[long_cpuid905])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc905_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid905/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 905 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid905]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc905_phy_pc_w))
                begin
                    if(good[long_cpuid905/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid905 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid905/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid905])
        end // if (done[905])

        if (done[906]) begin
            timeout[long_cpuid906] = 0;
            //check_bad_trap(spc906_phy_pc_w, 906, long_cpuid906);
            if(active_thread[long_cpuid906])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc906_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid906/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 906 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid906]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc906_phy_pc_w))
                begin
                    if(good[long_cpuid906/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid906 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid906/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid906])
        end // if (done[906])

        if (done[907]) begin
            timeout[long_cpuid907] = 0;
            //check_bad_trap(spc907_phy_pc_w, 907, long_cpuid907);
            if(active_thread[long_cpuid907])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc907_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid907/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 907 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid907]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc907_phy_pc_w))
                begin
                    if(good[long_cpuid907/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid907 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid907/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid907])
        end // if (done[907])

        if (done[908]) begin
            timeout[long_cpuid908] = 0;
            //check_bad_trap(spc908_phy_pc_w, 908, long_cpuid908);
            if(active_thread[long_cpuid908])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc908_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid908/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 908 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid908]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc908_phy_pc_w))
                begin
                    if(good[long_cpuid908/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid908 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid908/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid908])
        end // if (done[908])

        if (done[909]) begin
            timeout[long_cpuid909] = 0;
            //check_bad_trap(spc909_phy_pc_w, 909, long_cpuid909);
            if(active_thread[long_cpuid909])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc909_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid909/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 909 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid909]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc909_phy_pc_w))
                begin
                    if(good[long_cpuid909/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid909 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid909/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid909])
        end // if (done[909])

        if (done[910]) begin
            timeout[long_cpuid910] = 0;
            //check_bad_trap(spc910_phy_pc_w, 910, long_cpuid910);
            if(active_thread[long_cpuid910])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc910_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid910/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 910 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid910]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc910_phy_pc_w))
                begin
                    if(good[long_cpuid910/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid910 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid910/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid910])
        end // if (done[910])

        if (done[911]) begin
            timeout[long_cpuid911] = 0;
            //check_bad_trap(spc911_phy_pc_w, 911, long_cpuid911);
            if(active_thread[long_cpuid911])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc911_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid911/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 911 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid911]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc911_phy_pc_w))
                begin
                    if(good[long_cpuid911/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid911 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid911/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid911])
        end // if (done[911])

        if (done[912]) begin
            timeout[long_cpuid912] = 0;
            //check_bad_trap(spc912_phy_pc_w, 912, long_cpuid912);
            if(active_thread[long_cpuid912])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc912_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid912/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 912 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid912]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc912_phy_pc_w))
                begin
                    if(good[long_cpuid912/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid912 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid912/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid912])
        end // if (done[912])

        if (done[913]) begin
            timeout[long_cpuid913] = 0;
            //check_bad_trap(spc913_phy_pc_w, 913, long_cpuid913);
            if(active_thread[long_cpuid913])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc913_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid913/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 913 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid913]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc913_phy_pc_w))
                begin
                    if(good[long_cpuid913/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid913 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid913/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid913])
        end // if (done[913])

        if (done[914]) begin
            timeout[long_cpuid914] = 0;
            //check_bad_trap(spc914_phy_pc_w, 914, long_cpuid914);
            if(active_thread[long_cpuid914])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc914_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid914/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 914 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid914]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc914_phy_pc_w))
                begin
                    if(good[long_cpuid914/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid914 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid914/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid914])
        end // if (done[914])

        if (done[915]) begin
            timeout[long_cpuid915] = 0;
            //check_bad_trap(spc915_phy_pc_w, 915, long_cpuid915);
            if(active_thread[long_cpuid915])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc915_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid915/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 915 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid915]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc915_phy_pc_w))
                begin
                    if(good[long_cpuid915/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid915 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid915/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid915])
        end // if (done[915])

        if (done[916]) begin
            timeout[long_cpuid916] = 0;
            //check_bad_trap(spc916_phy_pc_w, 916, long_cpuid916);
            if(active_thread[long_cpuid916])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc916_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid916/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 916 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid916]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc916_phy_pc_w))
                begin
                    if(good[long_cpuid916/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid916 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid916/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid916])
        end // if (done[916])

        if (done[917]) begin
            timeout[long_cpuid917] = 0;
            //check_bad_trap(spc917_phy_pc_w, 917, long_cpuid917);
            if(active_thread[long_cpuid917])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc917_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid917/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 917 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid917]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc917_phy_pc_w))
                begin
                    if(good[long_cpuid917/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid917 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid917/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid917])
        end // if (done[917])

        if (done[918]) begin
            timeout[long_cpuid918] = 0;
            //check_bad_trap(spc918_phy_pc_w, 918, long_cpuid918);
            if(active_thread[long_cpuid918])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc918_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid918/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 918 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid918]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc918_phy_pc_w))
                begin
                    if(good[long_cpuid918/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid918 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid918/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid918])
        end // if (done[918])

        if (done[919]) begin
            timeout[long_cpuid919] = 0;
            //check_bad_trap(spc919_phy_pc_w, 919, long_cpuid919);
            if(active_thread[long_cpuid919])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc919_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid919/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 919 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid919]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc919_phy_pc_w))
                begin
                    if(good[long_cpuid919/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid919 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid919/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid919])
        end // if (done[919])

        if (done[920]) begin
            timeout[long_cpuid920] = 0;
            //check_bad_trap(spc920_phy_pc_w, 920, long_cpuid920);
            if(active_thread[long_cpuid920])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc920_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid920/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 920 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid920]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc920_phy_pc_w))
                begin
                    if(good[long_cpuid920/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid920 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid920/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid920])
        end // if (done[920])

        if (done[921]) begin
            timeout[long_cpuid921] = 0;
            //check_bad_trap(spc921_phy_pc_w, 921, long_cpuid921);
            if(active_thread[long_cpuid921])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc921_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid921/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 921 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid921]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc921_phy_pc_w))
                begin
                    if(good[long_cpuid921/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid921 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid921/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid921])
        end // if (done[921])

        if (done[922]) begin
            timeout[long_cpuid922] = 0;
            //check_bad_trap(spc922_phy_pc_w, 922, long_cpuid922);
            if(active_thread[long_cpuid922])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc922_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid922/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 922 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid922]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc922_phy_pc_w))
                begin
                    if(good[long_cpuid922/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid922 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid922/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid922])
        end // if (done[922])

        if (done[923]) begin
            timeout[long_cpuid923] = 0;
            //check_bad_trap(spc923_phy_pc_w, 923, long_cpuid923);
            if(active_thread[long_cpuid923])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc923_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid923/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 923 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid923]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc923_phy_pc_w))
                begin
                    if(good[long_cpuid923/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid923 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid923/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid923])
        end // if (done[923])

        if (done[924]) begin
            timeout[long_cpuid924] = 0;
            //check_bad_trap(spc924_phy_pc_w, 924, long_cpuid924);
            if(active_thread[long_cpuid924])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc924_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid924/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 924 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid924]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc924_phy_pc_w))
                begin
                    if(good[long_cpuid924/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid924 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid924/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid924])
        end // if (done[924])

        if (done[925]) begin
            timeout[long_cpuid925] = 0;
            //check_bad_trap(spc925_phy_pc_w, 925, long_cpuid925);
            if(active_thread[long_cpuid925])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc925_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid925/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 925 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid925]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc925_phy_pc_w))
                begin
                    if(good[long_cpuid925/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid925 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid925/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid925])
        end // if (done[925])

        if (done[926]) begin
            timeout[long_cpuid926] = 0;
            //check_bad_trap(spc926_phy_pc_w, 926, long_cpuid926);
            if(active_thread[long_cpuid926])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc926_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid926/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 926 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid926]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc926_phy_pc_w))
                begin
                    if(good[long_cpuid926/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid926 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid926/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid926])
        end // if (done[926])

        if (done[927]) begin
            timeout[long_cpuid927] = 0;
            //check_bad_trap(spc927_phy_pc_w, 927, long_cpuid927);
            if(active_thread[long_cpuid927])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc927_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid927/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 927 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid927]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc927_phy_pc_w))
                begin
                    if(good[long_cpuid927/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid927 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid927/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid927])
        end // if (done[927])

        if (done[928]) begin
            timeout[long_cpuid928] = 0;
            //check_bad_trap(spc928_phy_pc_w, 928, long_cpuid928);
            if(active_thread[long_cpuid928])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc928_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid928/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 928 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid928]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc928_phy_pc_w))
                begin
                    if(good[long_cpuid928/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid928 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid928/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid928])
        end // if (done[928])

        if (done[929]) begin
            timeout[long_cpuid929] = 0;
            //check_bad_trap(spc929_phy_pc_w, 929, long_cpuid929);
            if(active_thread[long_cpuid929])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc929_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid929/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 929 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid929]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc929_phy_pc_w))
                begin
                    if(good[long_cpuid929/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid929 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid929/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid929])
        end // if (done[929])

        if (done[930]) begin
            timeout[long_cpuid930] = 0;
            //check_bad_trap(spc930_phy_pc_w, 930, long_cpuid930);
            if(active_thread[long_cpuid930])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc930_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid930/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 930 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid930]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc930_phy_pc_w))
                begin
                    if(good[long_cpuid930/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid930 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid930/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid930])
        end // if (done[930])

        if (done[931]) begin
            timeout[long_cpuid931] = 0;
            //check_bad_trap(spc931_phy_pc_w, 931, long_cpuid931);
            if(active_thread[long_cpuid931])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc931_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid931/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 931 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid931]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc931_phy_pc_w))
                begin
                    if(good[long_cpuid931/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid931 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid931/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid931])
        end // if (done[931])

        if (done[932]) begin
            timeout[long_cpuid932] = 0;
            //check_bad_trap(spc932_phy_pc_w, 932, long_cpuid932);
            if(active_thread[long_cpuid932])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc932_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid932/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 932 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid932]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc932_phy_pc_w))
                begin
                    if(good[long_cpuid932/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid932 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid932/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid932])
        end // if (done[932])

        if (done[933]) begin
            timeout[long_cpuid933] = 0;
            //check_bad_trap(spc933_phy_pc_w, 933, long_cpuid933);
            if(active_thread[long_cpuid933])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc933_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid933/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 933 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid933]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc933_phy_pc_w))
                begin
                    if(good[long_cpuid933/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid933 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid933/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid933])
        end // if (done[933])

        if (done[934]) begin
            timeout[long_cpuid934] = 0;
            //check_bad_trap(spc934_phy_pc_w, 934, long_cpuid934);
            if(active_thread[long_cpuid934])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc934_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid934/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 934 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid934]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc934_phy_pc_w))
                begin
                    if(good[long_cpuid934/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid934 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid934/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid934])
        end // if (done[934])

        if (done[935]) begin
            timeout[long_cpuid935] = 0;
            //check_bad_trap(spc935_phy_pc_w, 935, long_cpuid935);
            if(active_thread[long_cpuid935])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc935_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid935/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 935 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid935]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc935_phy_pc_w))
                begin
                    if(good[long_cpuid935/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid935 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid935/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid935])
        end // if (done[935])

        if (done[936]) begin
            timeout[long_cpuid936] = 0;
            //check_bad_trap(spc936_phy_pc_w, 936, long_cpuid936);
            if(active_thread[long_cpuid936])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc936_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid936/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 936 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid936]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc936_phy_pc_w))
                begin
                    if(good[long_cpuid936/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid936 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid936/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid936])
        end // if (done[936])

        if (done[937]) begin
            timeout[long_cpuid937] = 0;
            //check_bad_trap(spc937_phy_pc_w, 937, long_cpuid937);
            if(active_thread[long_cpuid937])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc937_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid937/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 937 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid937]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc937_phy_pc_w))
                begin
                    if(good[long_cpuid937/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid937 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid937/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid937])
        end // if (done[937])

        if (done[938]) begin
            timeout[long_cpuid938] = 0;
            //check_bad_trap(spc938_phy_pc_w, 938, long_cpuid938);
            if(active_thread[long_cpuid938])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc938_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid938/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 938 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid938]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc938_phy_pc_w))
                begin
                    if(good[long_cpuid938/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid938 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid938/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid938])
        end // if (done[938])

        if (done[939]) begin
            timeout[long_cpuid939] = 0;
            //check_bad_trap(spc939_phy_pc_w, 939, long_cpuid939);
            if(active_thread[long_cpuid939])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc939_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid939/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 939 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid939]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc939_phy_pc_w))
                begin
                    if(good[long_cpuid939/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid939 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid939/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid939])
        end // if (done[939])

        if (done[940]) begin
            timeout[long_cpuid940] = 0;
            //check_bad_trap(spc940_phy_pc_w, 940, long_cpuid940);
            if(active_thread[long_cpuid940])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc940_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid940/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 940 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid940]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc940_phy_pc_w))
                begin
                    if(good[long_cpuid940/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid940 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid940/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid940])
        end // if (done[940])

        if (done[941]) begin
            timeout[long_cpuid941] = 0;
            //check_bad_trap(spc941_phy_pc_w, 941, long_cpuid941);
            if(active_thread[long_cpuid941])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc941_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid941/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 941 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid941]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc941_phy_pc_w))
                begin
                    if(good[long_cpuid941/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid941 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid941/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid941])
        end // if (done[941])

        if (done[942]) begin
            timeout[long_cpuid942] = 0;
            //check_bad_trap(spc942_phy_pc_w, 942, long_cpuid942);
            if(active_thread[long_cpuid942])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc942_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid942/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 942 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid942]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc942_phy_pc_w))
                begin
                    if(good[long_cpuid942/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid942 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid942/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid942])
        end // if (done[942])

        if (done[943]) begin
            timeout[long_cpuid943] = 0;
            //check_bad_trap(spc943_phy_pc_w, 943, long_cpuid943);
            if(active_thread[long_cpuid943])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc943_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid943/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 943 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid943]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc943_phy_pc_w))
                begin
                    if(good[long_cpuid943/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid943 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid943/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid943])
        end // if (done[943])

        if (done[944]) begin
            timeout[long_cpuid944] = 0;
            //check_bad_trap(spc944_phy_pc_w, 944, long_cpuid944);
            if(active_thread[long_cpuid944])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc944_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid944/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 944 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid944]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc944_phy_pc_w))
                begin
                    if(good[long_cpuid944/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid944 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid944/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid944])
        end // if (done[944])

        if (done[945]) begin
            timeout[long_cpuid945] = 0;
            //check_bad_trap(spc945_phy_pc_w, 945, long_cpuid945);
            if(active_thread[long_cpuid945])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc945_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid945/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 945 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid945]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc945_phy_pc_w))
                begin
                    if(good[long_cpuid945/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid945 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid945/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid945])
        end // if (done[945])

        if (done[946]) begin
            timeout[long_cpuid946] = 0;
            //check_bad_trap(spc946_phy_pc_w, 946, long_cpuid946);
            if(active_thread[long_cpuid946])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc946_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid946/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 946 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid946]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc946_phy_pc_w))
                begin
                    if(good[long_cpuid946/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid946 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid946/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid946])
        end // if (done[946])

        if (done[947]) begin
            timeout[long_cpuid947] = 0;
            //check_bad_trap(spc947_phy_pc_w, 947, long_cpuid947);
            if(active_thread[long_cpuid947])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc947_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid947/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 947 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid947]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc947_phy_pc_w))
                begin
                    if(good[long_cpuid947/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid947 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid947/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid947])
        end // if (done[947])

        if (done[948]) begin
            timeout[long_cpuid948] = 0;
            //check_bad_trap(spc948_phy_pc_w, 948, long_cpuid948);
            if(active_thread[long_cpuid948])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc948_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid948/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 948 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid948]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc948_phy_pc_w))
                begin
                    if(good[long_cpuid948/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid948 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid948/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid948])
        end // if (done[948])

        if (done[949]) begin
            timeout[long_cpuid949] = 0;
            //check_bad_trap(spc949_phy_pc_w, 949, long_cpuid949);
            if(active_thread[long_cpuid949])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc949_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid949/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 949 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid949]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc949_phy_pc_w))
                begin
                    if(good[long_cpuid949/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid949 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid949/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid949])
        end // if (done[949])

        if (done[950]) begin
            timeout[long_cpuid950] = 0;
            //check_bad_trap(spc950_phy_pc_w, 950, long_cpuid950);
            if(active_thread[long_cpuid950])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc950_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid950/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 950 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid950]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc950_phy_pc_w))
                begin
                    if(good[long_cpuid950/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid950 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid950/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid950])
        end // if (done[950])

        if (done[951]) begin
            timeout[long_cpuid951] = 0;
            //check_bad_trap(spc951_phy_pc_w, 951, long_cpuid951);
            if(active_thread[long_cpuid951])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc951_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid951/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 951 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid951]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc951_phy_pc_w))
                begin
                    if(good[long_cpuid951/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid951 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid951/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid951])
        end // if (done[951])

        if (done[952]) begin
            timeout[long_cpuid952] = 0;
            //check_bad_trap(spc952_phy_pc_w, 952, long_cpuid952);
            if(active_thread[long_cpuid952])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc952_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid952/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 952 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid952]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc952_phy_pc_w))
                begin
                    if(good[long_cpuid952/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid952 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid952/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid952])
        end // if (done[952])

        if (done[953]) begin
            timeout[long_cpuid953] = 0;
            //check_bad_trap(spc953_phy_pc_w, 953, long_cpuid953);
            if(active_thread[long_cpuid953])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc953_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid953/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 953 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid953]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc953_phy_pc_w))
                begin
                    if(good[long_cpuid953/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid953 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid953/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid953])
        end // if (done[953])

        if (done[954]) begin
            timeout[long_cpuid954] = 0;
            //check_bad_trap(spc954_phy_pc_w, 954, long_cpuid954);
            if(active_thread[long_cpuid954])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc954_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid954/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 954 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid954]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc954_phy_pc_w))
                begin
                    if(good[long_cpuid954/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid954 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid954/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid954])
        end // if (done[954])

        if (done[955]) begin
            timeout[long_cpuid955] = 0;
            //check_bad_trap(spc955_phy_pc_w, 955, long_cpuid955);
            if(active_thread[long_cpuid955])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc955_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid955/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 955 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid955]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc955_phy_pc_w))
                begin
                    if(good[long_cpuid955/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid955 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid955/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid955])
        end // if (done[955])

        if (done[956]) begin
            timeout[long_cpuid956] = 0;
            //check_bad_trap(spc956_phy_pc_w, 956, long_cpuid956);
            if(active_thread[long_cpuid956])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc956_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid956/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 956 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid956]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc956_phy_pc_w))
                begin
                    if(good[long_cpuid956/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid956 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid956/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid956])
        end // if (done[956])

        if (done[957]) begin
            timeout[long_cpuid957] = 0;
            //check_bad_trap(spc957_phy_pc_w, 957, long_cpuid957);
            if(active_thread[long_cpuid957])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc957_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid957/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 957 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid957]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc957_phy_pc_w))
                begin
                    if(good[long_cpuid957/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid957 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid957/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid957])
        end // if (done[957])

        if (done[958]) begin
            timeout[long_cpuid958] = 0;
            //check_bad_trap(spc958_phy_pc_w, 958, long_cpuid958);
            if(active_thread[long_cpuid958])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc958_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid958/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 958 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid958]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc958_phy_pc_w))
                begin
                    if(good[long_cpuid958/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid958 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid958/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid958])
        end // if (done[958])

        if (done[959]) begin
            timeout[long_cpuid959] = 0;
            //check_bad_trap(spc959_phy_pc_w, 959, long_cpuid959);
            if(active_thread[long_cpuid959])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc959_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid959/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 959 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid959]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc959_phy_pc_w))
                begin
                    if(good[long_cpuid959/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid959 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid959/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid959])
        end // if (done[959])

        if (done[960]) begin
            timeout[long_cpuid960] = 0;
            //check_bad_trap(spc960_phy_pc_w, 960, long_cpuid960);
            if(active_thread[long_cpuid960])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc960_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid960/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 960 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid960]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc960_phy_pc_w))
                begin
                    if(good[long_cpuid960/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid960 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid960/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid960])
        end // if (done[960])

        if (done[961]) begin
            timeout[long_cpuid961] = 0;
            //check_bad_trap(spc961_phy_pc_w, 961, long_cpuid961);
            if(active_thread[long_cpuid961])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc961_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid961/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 961 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid961]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc961_phy_pc_w))
                begin
                    if(good[long_cpuid961/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid961 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid961/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid961])
        end // if (done[961])

        if (done[962]) begin
            timeout[long_cpuid962] = 0;
            //check_bad_trap(spc962_phy_pc_w, 962, long_cpuid962);
            if(active_thread[long_cpuid962])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc962_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid962/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 962 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid962]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc962_phy_pc_w))
                begin
                    if(good[long_cpuid962/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid962 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid962/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid962])
        end // if (done[962])

        if (done[963]) begin
            timeout[long_cpuid963] = 0;
            //check_bad_trap(spc963_phy_pc_w, 963, long_cpuid963);
            if(active_thread[long_cpuid963])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc963_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid963/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 963 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid963]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc963_phy_pc_w))
                begin
                    if(good[long_cpuid963/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid963 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid963/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid963])
        end // if (done[963])

        if (done[964]) begin
            timeout[long_cpuid964] = 0;
            //check_bad_trap(spc964_phy_pc_w, 964, long_cpuid964);
            if(active_thread[long_cpuid964])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc964_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid964/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 964 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid964]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc964_phy_pc_w))
                begin
                    if(good[long_cpuid964/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid964 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid964/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid964])
        end // if (done[964])

        if (done[965]) begin
            timeout[long_cpuid965] = 0;
            //check_bad_trap(spc965_phy_pc_w, 965, long_cpuid965);
            if(active_thread[long_cpuid965])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc965_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid965/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 965 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid965]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc965_phy_pc_w))
                begin
                    if(good[long_cpuid965/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid965 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid965/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid965])
        end // if (done[965])

        if (done[966]) begin
            timeout[long_cpuid966] = 0;
            //check_bad_trap(spc966_phy_pc_w, 966, long_cpuid966);
            if(active_thread[long_cpuid966])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc966_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid966/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 966 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid966]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc966_phy_pc_w))
                begin
                    if(good[long_cpuid966/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid966 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid966/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid966])
        end // if (done[966])

        if (done[967]) begin
            timeout[long_cpuid967] = 0;
            //check_bad_trap(spc967_phy_pc_w, 967, long_cpuid967);
            if(active_thread[long_cpuid967])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc967_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid967/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 967 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid967]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc967_phy_pc_w))
                begin
                    if(good[long_cpuid967/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid967 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid967/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid967])
        end // if (done[967])

        if (done[968]) begin
            timeout[long_cpuid968] = 0;
            //check_bad_trap(spc968_phy_pc_w, 968, long_cpuid968);
            if(active_thread[long_cpuid968])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc968_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid968/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 968 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid968]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc968_phy_pc_w))
                begin
                    if(good[long_cpuid968/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid968 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid968/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid968])
        end // if (done[968])

        if (done[969]) begin
            timeout[long_cpuid969] = 0;
            //check_bad_trap(spc969_phy_pc_w, 969, long_cpuid969);
            if(active_thread[long_cpuid969])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc969_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid969/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 969 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid969]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc969_phy_pc_w))
                begin
                    if(good[long_cpuid969/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid969 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid969/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid969])
        end // if (done[969])

        if (done[970]) begin
            timeout[long_cpuid970] = 0;
            //check_bad_trap(spc970_phy_pc_w, 970, long_cpuid970);
            if(active_thread[long_cpuid970])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc970_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid970/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 970 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid970]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc970_phy_pc_w))
                begin
                    if(good[long_cpuid970/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid970 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid970/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid970])
        end // if (done[970])

        if (done[971]) begin
            timeout[long_cpuid971] = 0;
            //check_bad_trap(spc971_phy_pc_w, 971, long_cpuid971);
            if(active_thread[long_cpuid971])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc971_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid971/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 971 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid971]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc971_phy_pc_w))
                begin
                    if(good[long_cpuid971/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid971 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid971/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid971])
        end // if (done[971])

        if (done[972]) begin
            timeout[long_cpuid972] = 0;
            //check_bad_trap(spc972_phy_pc_w, 972, long_cpuid972);
            if(active_thread[long_cpuid972])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc972_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid972/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 972 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid972]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc972_phy_pc_w))
                begin
                    if(good[long_cpuid972/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid972 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid972/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid972])
        end // if (done[972])

        if (done[973]) begin
            timeout[long_cpuid973] = 0;
            //check_bad_trap(spc973_phy_pc_w, 973, long_cpuid973);
            if(active_thread[long_cpuid973])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc973_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid973/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 973 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid973]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc973_phy_pc_w))
                begin
                    if(good[long_cpuid973/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid973 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid973/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid973])
        end // if (done[973])

        if (done[974]) begin
            timeout[long_cpuid974] = 0;
            //check_bad_trap(spc974_phy_pc_w, 974, long_cpuid974);
            if(active_thread[long_cpuid974])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc974_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid974/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 974 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid974]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc974_phy_pc_w))
                begin
                    if(good[long_cpuid974/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid974 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid974/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid974])
        end // if (done[974])

        if (done[975]) begin
            timeout[long_cpuid975] = 0;
            //check_bad_trap(spc975_phy_pc_w, 975, long_cpuid975);
            if(active_thread[long_cpuid975])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc975_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid975/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 975 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid975]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc975_phy_pc_w))
                begin
                    if(good[long_cpuid975/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid975 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid975/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid975])
        end // if (done[975])

        if (done[976]) begin
            timeout[long_cpuid976] = 0;
            //check_bad_trap(spc976_phy_pc_w, 976, long_cpuid976);
            if(active_thread[long_cpuid976])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc976_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid976/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 976 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid976]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc976_phy_pc_w))
                begin
                    if(good[long_cpuid976/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid976 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid976/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid976])
        end // if (done[976])

        if (done[977]) begin
            timeout[long_cpuid977] = 0;
            //check_bad_trap(spc977_phy_pc_w, 977, long_cpuid977);
            if(active_thread[long_cpuid977])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc977_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid977/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 977 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid977]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc977_phy_pc_w))
                begin
                    if(good[long_cpuid977/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid977 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid977/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid977])
        end // if (done[977])

        if (done[978]) begin
            timeout[long_cpuid978] = 0;
            //check_bad_trap(spc978_phy_pc_w, 978, long_cpuid978);
            if(active_thread[long_cpuid978])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc978_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid978/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 978 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid978]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc978_phy_pc_w))
                begin
                    if(good[long_cpuid978/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid978 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid978/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid978])
        end // if (done[978])

        if (done[979]) begin
            timeout[long_cpuid979] = 0;
            //check_bad_trap(spc979_phy_pc_w, 979, long_cpuid979);
            if(active_thread[long_cpuid979])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc979_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid979/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 979 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid979]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc979_phy_pc_w))
                begin
                    if(good[long_cpuid979/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid979 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid979/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid979])
        end // if (done[979])

        if (done[980]) begin
            timeout[long_cpuid980] = 0;
            //check_bad_trap(spc980_phy_pc_w, 980, long_cpuid980);
            if(active_thread[long_cpuid980])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc980_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid980/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 980 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid980]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc980_phy_pc_w))
                begin
                    if(good[long_cpuid980/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid980 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid980/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid980])
        end // if (done[980])

        if (done[981]) begin
            timeout[long_cpuid981] = 0;
            //check_bad_trap(spc981_phy_pc_w, 981, long_cpuid981);
            if(active_thread[long_cpuid981])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc981_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid981/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 981 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid981]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc981_phy_pc_w))
                begin
                    if(good[long_cpuid981/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid981 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid981/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid981])
        end // if (done[981])

        if (done[982]) begin
            timeout[long_cpuid982] = 0;
            //check_bad_trap(spc982_phy_pc_w, 982, long_cpuid982);
            if(active_thread[long_cpuid982])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc982_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid982/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 982 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid982]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc982_phy_pc_w))
                begin
                    if(good[long_cpuid982/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid982 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid982/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid982])
        end // if (done[982])

        if (done[983]) begin
            timeout[long_cpuid983] = 0;
            //check_bad_trap(spc983_phy_pc_w, 983, long_cpuid983);
            if(active_thread[long_cpuid983])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc983_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid983/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 983 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid983]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc983_phy_pc_w))
                begin
                    if(good[long_cpuid983/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid983 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid983/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid983])
        end // if (done[983])

        if (done[984]) begin
            timeout[long_cpuid984] = 0;
            //check_bad_trap(spc984_phy_pc_w, 984, long_cpuid984);
            if(active_thread[long_cpuid984])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc984_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid984/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 984 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid984]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc984_phy_pc_w))
                begin
                    if(good[long_cpuid984/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid984 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid984/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid984])
        end // if (done[984])

        if (done[985]) begin
            timeout[long_cpuid985] = 0;
            //check_bad_trap(spc985_phy_pc_w, 985, long_cpuid985);
            if(active_thread[long_cpuid985])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc985_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid985/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 985 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid985]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc985_phy_pc_w))
                begin
                    if(good[long_cpuid985/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid985 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid985/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid985])
        end // if (done[985])

        if (done[986]) begin
            timeout[long_cpuid986] = 0;
            //check_bad_trap(spc986_phy_pc_w, 986, long_cpuid986);
            if(active_thread[long_cpuid986])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc986_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid986/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 986 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid986]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc986_phy_pc_w))
                begin
                    if(good[long_cpuid986/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid986 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid986/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid986])
        end // if (done[986])

        if (done[987]) begin
            timeout[long_cpuid987] = 0;
            //check_bad_trap(spc987_phy_pc_w, 987, long_cpuid987);
            if(active_thread[long_cpuid987])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc987_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid987/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 987 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid987]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc987_phy_pc_w))
                begin
                    if(good[long_cpuid987/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid987 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid987/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid987])
        end // if (done[987])

        if (done[988]) begin
            timeout[long_cpuid988] = 0;
            //check_bad_trap(spc988_phy_pc_w, 988, long_cpuid988);
            if(active_thread[long_cpuid988])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc988_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid988/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 988 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid988]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc988_phy_pc_w))
                begin
                    if(good[long_cpuid988/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid988 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid988/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid988])
        end // if (done[988])

        if (done[989]) begin
            timeout[long_cpuid989] = 0;
            //check_bad_trap(spc989_phy_pc_w, 989, long_cpuid989);
            if(active_thread[long_cpuid989])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc989_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid989/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 989 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid989]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc989_phy_pc_w))
                begin
                    if(good[long_cpuid989/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid989 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid989/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid989])
        end // if (done[989])

        if (done[990]) begin
            timeout[long_cpuid990] = 0;
            //check_bad_trap(spc990_phy_pc_w, 990, long_cpuid990);
            if(active_thread[long_cpuid990])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc990_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid990/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 990 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid990]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc990_phy_pc_w))
                begin
                    if(good[long_cpuid990/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid990 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid990/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid990])
        end // if (done[990])

        if (done[991]) begin
            timeout[long_cpuid991] = 0;
            //check_bad_trap(spc991_phy_pc_w, 991, long_cpuid991);
            if(active_thread[long_cpuid991])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc991_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid991/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 991 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid991]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc991_phy_pc_w))
                begin
                    if(good[long_cpuid991/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid991 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid991/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid991])
        end // if (done[991])

        if (done[992]) begin
            timeout[long_cpuid992] = 0;
            //check_bad_trap(spc992_phy_pc_w, 992, long_cpuid992);
            if(active_thread[long_cpuid992])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc992_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid992/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 992 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid992]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc992_phy_pc_w))
                begin
                    if(good[long_cpuid992/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid992 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid992/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid992])
        end // if (done[992])

        if (done[993]) begin
            timeout[long_cpuid993] = 0;
            //check_bad_trap(spc993_phy_pc_w, 993, long_cpuid993);
            if(active_thread[long_cpuid993])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc993_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid993/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 993 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid993]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc993_phy_pc_w))
                begin
                    if(good[long_cpuid993/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid993 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid993/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid993])
        end // if (done[993])

        if (done[994]) begin
            timeout[long_cpuid994] = 0;
            //check_bad_trap(spc994_phy_pc_w, 994, long_cpuid994);
            if(active_thread[long_cpuid994])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc994_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid994/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 994 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid994]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc994_phy_pc_w))
                begin
                    if(good[long_cpuid994/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid994 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid994/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid994])
        end // if (done[994])

        if (done[995]) begin
            timeout[long_cpuid995] = 0;
            //check_bad_trap(spc995_phy_pc_w, 995, long_cpuid995);
            if(active_thread[long_cpuid995])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc995_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid995/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 995 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid995]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc995_phy_pc_w))
                begin
                    if(good[long_cpuid995/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid995 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid995/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid995])
        end // if (done[995])

        if (done[996]) begin
            timeout[long_cpuid996] = 0;
            //check_bad_trap(spc996_phy_pc_w, 996, long_cpuid996);
            if(active_thread[long_cpuid996])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc996_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid996/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 996 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid996]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc996_phy_pc_w))
                begin
                    if(good[long_cpuid996/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid996 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid996/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid996])
        end // if (done[996])

        if (done[997]) begin
            timeout[long_cpuid997] = 0;
            //check_bad_trap(spc997_phy_pc_w, 997, long_cpuid997);
            if(active_thread[long_cpuid997])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc997_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid997/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 997 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid997]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc997_phy_pc_w))
                begin
                    if(good[long_cpuid997/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid997 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid997/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid997])
        end // if (done[997])

        if (done[998]) begin
            timeout[long_cpuid998] = 0;
            //check_bad_trap(spc998_phy_pc_w, 998, long_cpuid998);
            if(active_thread[long_cpuid998])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc998_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid998/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 998 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid998]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc998_phy_pc_w))
                begin
                    if(good[long_cpuid998/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid998 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid998/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid998])
        end // if (done[998])

        if (done[999]) begin
            timeout[long_cpuid999] = 0;
            //check_bad_trap(spc999_phy_pc_w, 999, long_cpuid999);
            if(active_thread[long_cpuid999])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc999_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid999/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 999 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid999]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc999_phy_pc_w))
                begin
                    if(good[long_cpuid999/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid999 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid999/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid999])
        end // if (done[999])

        if (done[1000]) begin
            timeout[long_cpuid1000] = 0;
            //check_bad_trap(spc1000_phy_pc_w, 1000, long_cpuid1000);
            if(active_thread[long_cpuid1000])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc1000_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid1000/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 1000 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid1000]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc1000_phy_pc_w))
                begin
                    if(good[long_cpuid1000/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid1000 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid1000/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid1000])
        end // if (done[1000])

        if (done[1001]) begin
            timeout[long_cpuid1001] = 0;
            //check_bad_trap(spc1001_phy_pc_w, 1001, long_cpuid1001);
            if(active_thread[long_cpuid1001])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc1001_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid1001/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 1001 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid1001]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc1001_phy_pc_w))
                begin
                    if(good[long_cpuid1001/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid1001 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid1001/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid1001])
        end // if (done[1001])

        if (done[1002]) begin
            timeout[long_cpuid1002] = 0;
            //check_bad_trap(spc1002_phy_pc_w, 1002, long_cpuid1002);
            if(active_thread[long_cpuid1002])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc1002_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid1002/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 1002 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid1002]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc1002_phy_pc_w))
                begin
                    if(good[long_cpuid1002/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid1002 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid1002/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid1002])
        end // if (done[1002])

        if (done[1003]) begin
            timeout[long_cpuid1003] = 0;
            //check_bad_trap(spc1003_phy_pc_w, 1003, long_cpuid1003);
            if(active_thread[long_cpuid1003])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc1003_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid1003/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 1003 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid1003]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc1003_phy_pc_w))
                begin
                    if(good[long_cpuid1003/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid1003 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid1003/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid1003])
        end // if (done[1003])

        if (done[1004]) begin
            timeout[long_cpuid1004] = 0;
            //check_bad_trap(spc1004_phy_pc_w, 1004, long_cpuid1004);
            if(active_thread[long_cpuid1004])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc1004_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid1004/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 1004 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid1004]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc1004_phy_pc_w))
                begin
                    if(good[long_cpuid1004/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid1004 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid1004/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid1004])
        end // if (done[1004])

        if (done[1005]) begin
            timeout[long_cpuid1005] = 0;
            //check_bad_trap(spc1005_phy_pc_w, 1005, long_cpuid1005);
            if(active_thread[long_cpuid1005])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc1005_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid1005/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 1005 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid1005]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc1005_phy_pc_w))
                begin
                    if(good[long_cpuid1005/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid1005 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid1005/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid1005])
        end // if (done[1005])

        if (done[1006]) begin
            timeout[long_cpuid1006] = 0;
            //check_bad_trap(spc1006_phy_pc_w, 1006, long_cpuid1006);
            if(active_thread[long_cpuid1006])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc1006_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid1006/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 1006 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid1006]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc1006_phy_pc_w))
                begin
                    if(good[long_cpuid1006/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid1006 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid1006/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid1006])
        end // if (done[1006])

        if (done[1007]) begin
            timeout[long_cpuid1007] = 0;
            //check_bad_trap(spc1007_phy_pc_w, 1007, long_cpuid1007);
            if(active_thread[long_cpuid1007])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc1007_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid1007/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 1007 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid1007]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc1007_phy_pc_w))
                begin
                    if(good[long_cpuid1007/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid1007 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid1007/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid1007])
        end // if (done[1007])

        if (done[1008]) begin
            timeout[long_cpuid1008] = 0;
            //check_bad_trap(spc1008_phy_pc_w, 1008, long_cpuid1008);
            if(active_thread[long_cpuid1008])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc1008_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid1008/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 1008 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid1008]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc1008_phy_pc_w))
                begin
                    if(good[long_cpuid1008/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid1008 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid1008/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid1008])
        end // if (done[1008])

        if (done[1009]) begin
            timeout[long_cpuid1009] = 0;
            //check_bad_trap(spc1009_phy_pc_w, 1009, long_cpuid1009);
            if(active_thread[long_cpuid1009])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc1009_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid1009/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 1009 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid1009]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc1009_phy_pc_w))
                begin
                    if(good[long_cpuid1009/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid1009 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid1009/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid1009])
        end // if (done[1009])

        if (done[1010]) begin
            timeout[long_cpuid1010] = 0;
            //check_bad_trap(spc1010_phy_pc_w, 1010, long_cpuid1010);
            if(active_thread[long_cpuid1010])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc1010_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid1010/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 1010 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid1010]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc1010_phy_pc_w))
                begin
                    if(good[long_cpuid1010/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid1010 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid1010/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid1010])
        end // if (done[1010])

        if (done[1011]) begin
            timeout[long_cpuid1011] = 0;
            //check_bad_trap(spc1011_phy_pc_w, 1011, long_cpuid1011);
            if(active_thread[long_cpuid1011])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc1011_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid1011/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 1011 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid1011]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc1011_phy_pc_w))
                begin
                    if(good[long_cpuid1011/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid1011 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid1011/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid1011])
        end // if (done[1011])

        if (done[1012]) begin
            timeout[long_cpuid1012] = 0;
            //check_bad_trap(spc1012_phy_pc_w, 1012, long_cpuid1012);
            if(active_thread[long_cpuid1012])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc1012_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid1012/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 1012 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid1012]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc1012_phy_pc_w))
                begin
                    if(good[long_cpuid1012/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid1012 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid1012/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid1012])
        end // if (done[1012])

        if (done[1013]) begin
            timeout[long_cpuid1013] = 0;
            //check_bad_trap(spc1013_phy_pc_w, 1013, long_cpuid1013);
            if(active_thread[long_cpuid1013])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc1013_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid1013/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 1013 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid1013]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc1013_phy_pc_w))
                begin
                    if(good[long_cpuid1013/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid1013 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid1013/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid1013])
        end // if (done[1013])

        if (done[1014]) begin
            timeout[long_cpuid1014] = 0;
            //check_bad_trap(spc1014_phy_pc_w, 1014, long_cpuid1014);
            if(active_thread[long_cpuid1014])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc1014_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid1014/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 1014 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid1014]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc1014_phy_pc_w))
                begin
                    if(good[long_cpuid1014/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid1014 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid1014/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid1014])
        end // if (done[1014])

        if (done[1015]) begin
            timeout[long_cpuid1015] = 0;
            //check_bad_trap(spc1015_phy_pc_w, 1015, long_cpuid1015);
            if(active_thread[long_cpuid1015])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc1015_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid1015/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 1015 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid1015]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc1015_phy_pc_w))
                begin
                    if(good[long_cpuid1015/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid1015 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid1015/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid1015])
        end // if (done[1015])

        if (done[1016]) begin
            timeout[long_cpuid1016] = 0;
            //check_bad_trap(spc1016_phy_pc_w, 1016, long_cpuid1016);
            if(active_thread[long_cpuid1016])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc1016_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid1016/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 1016 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid1016]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc1016_phy_pc_w))
                begin
                    if(good[long_cpuid1016/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid1016 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid1016/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid1016])
        end // if (done[1016])

        if (done[1017]) begin
            timeout[long_cpuid1017] = 0;
            //check_bad_trap(spc1017_phy_pc_w, 1017, long_cpuid1017);
            if(active_thread[long_cpuid1017])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc1017_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid1017/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 1017 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid1017]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc1017_phy_pc_w))
                begin
                    if(good[long_cpuid1017/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid1017 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid1017/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid1017])
        end // if (done[1017])

        if (done[1018]) begin
            timeout[long_cpuid1018] = 0;
            //check_bad_trap(spc1018_phy_pc_w, 1018, long_cpuid1018);
            if(active_thread[long_cpuid1018])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc1018_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid1018/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 1018 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid1018]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc1018_phy_pc_w))
                begin
                    if(good[long_cpuid1018/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid1018 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid1018/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid1018])
        end // if (done[1018])

        if (done[1019]) begin
            timeout[long_cpuid1019] = 0;
            //check_bad_trap(spc1019_phy_pc_w, 1019, long_cpuid1019);
            if(active_thread[long_cpuid1019])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc1019_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid1019/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 1019 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid1019]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc1019_phy_pc_w))
                begin
                    if(good[long_cpuid1019/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid1019 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid1019/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid1019])
        end // if (done[1019])

        if (done[1020]) begin
            timeout[long_cpuid1020] = 0;
            //check_bad_trap(spc1020_phy_pc_w, 1020, long_cpuid1020);
            if(active_thread[long_cpuid1020])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc1020_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid1020/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 1020 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid1020]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc1020_phy_pc_w))
                begin
                    if(good[long_cpuid1020/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid1020 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid1020/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid1020])
        end // if (done[1020])

        if (done[1021]) begin
            timeout[long_cpuid1021] = 0;
            //check_bad_trap(spc1021_phy_pc_w, 1021, long_cpuid1021);
            if(active_thread[long_cpuid1021])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc1021_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid1021/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 1021 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid1021]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc1021_phy_pc_w))
                begin
                    if(good[long_cpuid1021/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid1021 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid1021/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid1021])
        end // if (done[1021])

        if (done[1022]) begin
            timeout[long_cpuid1022] = 0;
            //check_bad_trap(spc1022_phy_pc_w, 1022, long_cpuid1022);
            if(active_thread[long_cpuid1022])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc1022_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid1022/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 1022 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid1022]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc1022_phy_pc_w))
                begin
                    if(good[long_cpuid1022/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid1022 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid1022/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid1022])
        end // if (done[1022])

        if (done[1023]) begin
            timeout[long_cpuid1023] = 0;
            //check_bad_trap(spc1023_phy_pc_w, 1023, long_cpuid1023);
            if(active_thread[long_cpuid1023])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc1023_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid1023/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 1023 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid1023]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc1023_phy_pc_w))
                begin
                    if(good[long_cpuid1023/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid1023 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid1023/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid1023])
        end // if (done[1023])

        
        end
`ifdef INCLUDE_SAS_TASKS
        get_thread_status;
`endif
        set_diag_done(local_diag_done);
    end // if (rst_l)
end // always @ (posedge clk)

always @(posedge clk) begin
  if (!rst_l) begin
    good <= '0;
    hit_bad <= 1'b0;
  end else begin
    if (&good) begin
      $display("All threads hit good tap - PASS");
      $finish;
    end
    if (hit_bad) begin
      $display("A thread hit bad trap - FAIL");
      $error;
      $finish;
    end
  end
end

endmodule


