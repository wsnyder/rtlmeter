// Modified by Princeton University on June 9th, 2015
// ========== Copyright Header Begin ==========================================
//
// OpenSPARC T1 Processor File: iop.v
// Copyright (c) 2006 Sun Microsystems, Inc.  All Rights Reserved.
// DO NOT ALTER OR REMOVE COPYRIGHT NOTICES.
//
// The above named program is free software; you can redistribute it and/or
// modify it under the terms of the GNU General Public
// License version 2 as published by the Free Software Foundation.
//
// The above named program is distributed in the hope that it will be
// useful, but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
// General Public License for more details.
//
// You should have received a copy of the GNU General Public
// License along with this work; if not, write to the Free Software
// Foundation, Inc., 51 Franklin St, Fifth Floor, Boston, MA 02110-1301, USA.
//
// ========== Copyright Header End ============================================

`ifndef USE_TEST_TOP // useless for older TOPs

`include "define.tmp.h"
`include "piton_system.vh"
`include "jtag.vh"

module chip(
`ifndef PITON_CHIP_FPGA
   // IO cell configs
   input                                        slew,
   input                                        impsel1,
   input                                        impsel2,
`endif // endif PITON_CHIP_FPGA

`ifdef PITON_FPGA_CLKS_GEN
   input                                        clk_osc_p,
   input                                        clk_osc_n,
`else // ifndef PITON_FPGA_CLKS_GEN
   // Input clocks
   input                                        core_ref_clk,
   input                                        io_clk,
`endif // endif PITON_FPGA_CLKS_GEN

   // Resets
   // reset is assumed to be asynchronous
   input                                        rst_n,
`ifndef PITON_CHIP_FPGA
   input                                        pll_rst_n,

   // Chip-level clock enable
   input                                        clk_en,

   // PLL settings
   output                                       pll_lock,
   input                                        pll_bypass,
   input  [4:0]                                 pll_rangea,

   // Clock mux select (bypass PLL or not)
   // Double redundancy with pll_bypass
   input  [1:0]                                 clk_mux_sel,

   // JTAG
   input                                        jtag_clk,
   input                                        jtag_rst_l,
   input                                        jtag_modesel,
   input                                        jtag_datain,
   output                                       jtag_dataout,

   // Async FIFOs enable
   input                                        async_mux,

   // ORAM
   input                                        oram_on,
   input                                        oram_traffic_gen,
   input                                        oram_dummy_gen,
`else // ifdef PITON_CHIP_FPGA
   // Need to output this to chipset, since there will
   // be no passthru in the case of synthesizing chip on its own
   output                                       piton_prsnt_n,
   output                                       piton_ready_n,

   input                                        chipset_prsnt_n,

   output [7:0]                                 leds,
`endif // endif PITON_CHIP_FPGA

`ifndef PITON_NO_CHIP_BRIDGE
   // For FPGA implementations, we convert to differential and source synchronous
`ifdef PITON_CHIP_FPGA
   output                                      chip_intf_clk_p,
   output                                      chip_intf_clk_n,
   input                                       intf_chip_clk_p,
   input                                       intf_chip_clk_n,

   output [31:0]                               chip_intf_data_p,
   output [31:0]                               chip_intf_data_n,
   output [1:0]                                chip_intf_channel_p,
   output [1:0]                                chip_intf_channel_n,
   input  [2:0]                                chip_intf_credit_back_p,
   input  [2:0]                                chip_intf_credit_back_n,

   input  [31:0]                               intf_chip_data_p,
   input  [31:0]                               intf_chip_data_n,
   input  [1:0]                                intf_chip_channel_p,
   input  [1:0]                                intf_chip_channel_n,
   output [2:0]                                intf_chip_credit_back_p,
   output [2:0]                                intf_chip_credit_back_n
`else // ifndef PITON_CHIP_FPGA
   // Virtual channel credit-based off-chip interface
   input  [31:0]                                intf_chip_data,
   input  [1:0]                                 intf_chip_channel,
   output [2:0]                                 intf_chip_credit_back,

   output [31:0]                                chip_intf_data,
   output [1:0]                                 chip_intf_channel,
   input  [2:0]                                 chip_intf_credit_back
`endif // endif PITON_CHIP_FPGA
`else // ifdef PITON_NO_CHIP_BRIDGE
   output                                       processor_offchip_noc1_valid,
   output [`NOC_DATA_WIDTH-1:0]                 processor_offchip_noc1_data,
   input                                        processor_offchip_noc1_yummy,
   output                                       processor_offchip_noc2_valid,
   output [`NOC_DATA_WIDTH-1:0]                 processor_offchip_noc2_data,
   input                                        processor_offchip_noc2_yummy,
   output                                       processor_offchip_noc3_valid,
   output [`NOC_DATA_WIDTH-1:0]                 processor_offchip_noc3_data,
   input                                        processor_offchip_noc3_yummy,

   input                                        offchip_processor_noc1_valid,
   input  [`NOC_DATA_WIDTH-1:0]                 offchip_processor_noc1_data,
   output                                       offchip_processor_noc1_yummy,
   input                                        offchip_processor_noc2_valid,
   input  [`NOC_DATA_WIDTH-1:0]                 offchip_processor_noc2_data,
   output                                       offchip_processor_noc2_yummy,
   input                                        offchip_processor_noc3_valid,
   input  [`NOC_DATA_WIDTH-1:0]                 offchip_processor_noc3_data,
   output                                       offchip_processor_noc3_yummy
`endif // endif PITON_NO_CHIP_BRIDGE

`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    // Debug
,   input                                       ndmreset_i      // non-debug module reset
,   input   [`PITON_NUM_TILES-1:0]              debug_req_i     // async debug request
,   output  [`PITON_NUM_TILES-1:0]              unavailable_o   // communicate whether the hart is unavailable (e.g.: power down)
`endif // ifdef PITON_RV64_DEBUGUNIT

`ifdef PITON_RV64_CLINT
    // CLINT
,   input   [`PITON_NUM_TILES-1:0]              timer_irq_i     // Timer interrupts
,   input   [`PITON_NUM_TILES-1:0]              ipi_i           // software interrupt (a.k.a inter-process-interrupt)
`endif // ifdef PITON_RV64_CLINT

`ifdef PITON_RV64_PLIC
    // PLIC
,   input   [`PITON_NUM_TILES*2-1:0]            irq_i           // level sensitive IR lines, mip & sip (async)
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
);

// /home/gl/work/openpiton/piton/verif/env/manycore/devices_ariane.xml


   ///////////////////////
   // Type Declarations
   ///////////////////////

   // Need to define types for missing inputs and outputs
   // if synthesizing chip to fpga standalone
`ifdef PITON_CHIP_FPGA
   wire                                         slew;
   wire                                         impsel1;
   wire                                         impsel2;


   wire                                         pll_rst_n;

   wire                                         clk_en;

   wire                                         pll_lock;
   wire                                         pll_bypass;
   wire [4:0]                                   pll_rangea;

   wire [1:0]                                   clk_mux_sel;

   wire                                         jtag_clk;
   wire                                         jtag_rst_l;
   wire                                         jtag_modesel;
   wire                                         jtag_datain;
   wire                                         jtag_dataout;

   wire                                         async_mux;

   wire                                         oram_on;
   wire                                         oram_traffic_gen;
   wire                                         oram_dummy_gen;
`endif // endif PITON_CHIP_FPGA
   // Same for generating clocks
`ifdef PITON_FPGA_CLKS_GEN
   wire                                         core_ref_clk;

   wire                                         mmcm_locked;
`endif // endif PITON_FPGA_CLKS_GEN
   // Same for chip interface
`ifndef PITON_NO_CHIP_BRIDGE
`ifdef PITON_CHIP_FPGA
   wire                                         io_clk;

   wire [31:0]                                  intf_chip_data;
   wire [1:0]                                   intf_chip_channel;
   wire [2:0]                                   intf_chip_credit_back;

   wire [31:0]                                  chip_intf_data;
   wire [1:0]                                   chip_intf_channel;
   wire [2:0]                                   chip_intf_credit_back;
`endif // endif PITON_CHIP_FPGA
`endif // endif PITON_NO_CHIP_BRIDGE

   // OCI internal wires

   wire                                         core_ref_clk_inter;
   wire                                         io_clk_inter;
   wire                                         rst_n_inter;
   wire                                         pll_rst_n_inter;
   wire                                         clk_en_inter;
   wire                                         pll_lock_inter;
   wire                                         pll_bypass_inter;
   wire [4:0]                                   pll_rangea_inter;
   wire [1:0]                                   clk_mux_sel_inter;
   wire                                         jtag_clk_inter;
   wire                                         jtag_rst_l_inter;
   wire                                         jtag_rst_l_inter_sync;
   wire                                         jtag_modesel_inter;
   wire                                         jtag_datain_inter;
   wire                                         jtag_dataout_inter;
   wire                                         async_mux_inter;
   wire                                         oram_on_inter;
   wire                                         oram_traffic_gen_inter;
   wire                                         oram_dummy_gen_inter;
   wire [31:0]                              intf_chip_data_inter;
   wire [1:0]                                   intf_chip_channel_inter;
   wire [2:0]                                   intf_chip_credit_back_inter;
   wire [31:0]                                  chip_intf_data_inter;
   wire [1:0]                                   chip_intf_channel_inter;
   wire [2:0]                                   chip_intf_credit_back_inter;

   // Synchronized resets
   wire                                         rst_n_inter_sync;
   reg                                          rst_n_inter_sync_f;
   wire                                         io_clk_rst_n_inter_sync;
   reg                                          io_clk_rst_n_inter_sync_f;

   // PLL signals
   wire                                         core_ref_clk_inter_c;
   wire                                         core_ref_clk_inter_t;
   wire                                         clk_muxed;
   wire                                         pll_clk;

   // Buffered chip bridge inputs
   reg  [31:0]                                  intf_chip_data_inter_buf_f /* synthesis iob = true */;
   reg  [1:0]                                   intf_chip_channel_inter_buf_f /* synthesis iob = true */;
   reg  [2:0]                                   chip_intf_credit_back_inter_buf_f /* synthesis iob = true */;

   // Chip bridge val/rdy interface
   wire                                         chip_intf_noc1_valid;
   wire [`NOC_DATA_WIDTH-1:0]                   chip_intf_noc1_data;
   wire                                         chip_intf_noc1_rdy;
   wire                                         chip_intf_noc2_valid;
   wire [`NOC_DATA_WIDTH-1:0]                   chip_intf_noc2_data;
   wire                                         chip_intf_noc2_rdy;
   wire                                         chip_intf_noc3_valid;
   wire [`NOC_DATA_WIDTH-1:0]                   chip_intf_noc3_data;
   wire                                         chip_intf_noc3_rdy;

   wire                                         intf_chip_noc1_valid;
   wire [`NOC_DATA_WIDTH-1:0]                   intf_chip_noc1_data;
   wire                                         intf_chip_noc1_rdy;
   wire                                         intf_chip_noc2_valid;
   wire [`NOC_DATA_WIDTH-1:0]                   intf_chip_noc2_data;
   wire                                         intf_chip_noc2_rdy;
   wire                                         intf_chip_noc3_valid;
   wire [`NOC_DATA_WIDTH-1:0]                   intf_chip_noc3_data;
   wire                                         intf_chip_noc3_rdy;

`ifndef PITON_NO_CHIP_BRIDGE
   // Need to convert a chip bridge interface to these if PITON_NO_CHIP_BRIDGE
   // is not specified
   wire                                         processor_offchip_noc1_valid;
   wire [`NOC_DATA_WIDTH-1:0]                   processor_offchip_noc1_data;
   wire                                         processor_offchip_noc1_yummy;
   wire                                         processor_offchip_noc2_valid;
   wire [`NOC_DATA_WIDTH-1:0]                   processor_offchip_noc2_data;
   wire                                         processor_offchip_noc2_yummy;
   wire                                         processor_offchip_noc3_valid;
   wire [`NOC_DATA_WIDTH-1:0]                   processor_offchip_noc3_data;
   wire                                         processor_offchip_noc3_yummy;

   wire                                         offchip_processor_noc1_valid;
   wire [`NOC_DATA_WIDTH-1:0]                   offchip_processor_noc1_data;
   wire                                         offchip_processor_noc1_yummy;
   wire                                         offchip_processor_noc2_valid;
   wire [`NOC_DATA_WIDTH-1:0]                   offchip_processor_noc2_data;
   wire                                         offchip_processor_noc2_yummy;
   wire                                         offchip_processor_noc3_valid;
   wire [`NOC_DATA_WIDTH-1:0]                   offchip_processor_noc3_data;
   wire                                         offchip_processor_noc3_yummy;
`endif // endif PITON_NO_CHIP_BRIDGE

   // ORAM muxed outputs
   reg                                          proc_oram_yummy;
   reg                                          oram_proc_valid;
   reg  [`NOC_DATA_WIDTH-1:0]                   oram_proc_data;
   reg                                          offchip_oram_yummy;
   reg                                          oram_offchip_valid;
   reg  [`NOC_DATA_WIDTH-1:0]                   oram_offchip_data;

   // ORAM Signals
   wire                                         proc_oram_valid;
   wire [`NOC_DATA_WIDTH-1:0]                   proc_oram_data;
   wire                                         proc_oram_yummy_oram;
   wire                                         oram_proc_valid_oram;
   wire [`NOC_DATA_WIDTH-1:0]                   oram_proc_data_oram;
   wire                                         oram_proc_yummy;

   wire                                         offchip_oram_valid;
   wire [`NOC_DATA_WIDTH-1:0]                   offchip_oram_data;
   wire                                         offchip_oram_yummy_oram;
   wire                                         oram_offchip_valid_oram;
   wire [`NOC_DATA_WIDTH-1:0]                   oram_offchip_data_oram;
   wire                                         oram_offchip_yummy;

   // ORAM JTAG Signals
   wire                                         ctap_oram_clk_en;
   wire                                         ctap_oram_req_val;
   wire [`JTAG_ORAM_MISC_WIDTH-1:0]             ctap_oram_req_misc;
   wire [`JTAG_ORAM_DATA_WIDTH-1:0]             oram_ctap_res_data;
   // wire [`BIST_OP_WIDTH-1:0]                    ctap_oram_bist_command;
   // wire [`SRAM_WRAPPER_BUS_WIDTH-1:0]           ctap_oram_bist_data;
   // wire [`SRAM_WRAPPER_BUS_WIDTH-1:0]           oram_ctap_sram_data;

   // Merged JTAG outputs from tile
   wire                                         tiles_jtag_ucb_val;
   wire [`UCB_BUS_WIDTH-1:0]                    tiles_jtag_ucb_data;

   // Tiles JTAG interface
   wire                                         jtag_tiles_ucb_val;
   wire [`UCB_BUS_WIDTH-1:0]                    jtag_tiles_ucb_data;
   wire [127:0]                                 ctap_clk_en_inter; // trin TODO: parameterize this number (63)
   wire tile0_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile0_jtag_ucb_data;
wire tile16_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile16_jtag_ucb_data;
wire tile32_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile32_jtag_ucb_data;
wire tile48_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile48_jtag_ucb_data;
wire tile64_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile64_jtag_ucb_data;
wire tile80_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile80_jtag_ucb_data;
wire tile96_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile96_jtag_ucb_data;
wire tile112_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile112_jtag_ucb_data;
wire tile128_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile128_jtag_ucb_data;
wire tile144_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile144_jtag_ucb_data;
wire tile160_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile160_jtag_ucb_data;
wire tile176_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile176_jtag_ucb_data;
wire tile192_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile192_jtag_ucb_data;
wire tile208_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile208_jtag_ucb_data;
wire tile224_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile224_jtag_ucb_data;
wire tile240_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile240_jtag_ucb_data;
wire tile1_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile1_jtag_ucb_data;
wire tile17_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile17_jtag_ucb_data;
wire tile33_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile33_jtag_ucb_data;
wire tile49_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile49_jtag_ucb_data;
wire tile65_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile65_jtag_ucb_data;
wire tile81_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile81_jtag_ucb_data;
wire tile97_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile97_jtag_ucb_data;
wire tile113_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile113_jtag_ucb_data;
wire tile129_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile129_jtag_ucb_data;
wire tile145_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile145_jtag_ucb_data;
wire tile161_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile161_jtag_ucb_data;
wire tile177_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile177_jtag_ucb_data;
wire tile193_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile193_jtag_ucb_data;
wire tile209_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile209_jtag_ucb_data;
wire tile225_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile225_jtag_ucb_data;
wire tile241_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile241_jtag_ucb_data;
wire tile2_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile2_jtag_ucb_data;
wire tile18_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile18_jtag_ucb_data;
wire tile34_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile34_jtag_ucb_data;
wire tile50_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile50_jtag_ucb_data;
wire tile66_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile66_jtag_ucb_data;
wire tile82_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile82_jtag_ucb_data;
wire tile98_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile98_jtag_ucb_data;
wire tile114_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile114_jtag_ucb_data;
wire tile130_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile130_jtag_ucb_data;
wire tile146_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile146_jtag_ucb_data;
wire tile162_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile162_jtag_ucb_data;
wire tile178_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile178_jtag_ucb_data;
wire tile194_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile194_jtag_ucb_data;
wire tile210_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile210_jtag_ucb_data;
wire tile226_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile226_jtag_ucb_data;
wire tile242_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile242_jtag_ucb_data;
wire tile3_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile3_jtag_ucb_data;
wire tile19_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile19_jtag_ucb_data;
wire tile35_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile35_jtag_ucb_data;
wire tile51_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile51_jtag_ucb_data;
wire tile67_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile67_jtag_ucb_data;
wire tile83_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile83_jtag_ucb_data;
wire tile99_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile99_jtag_ucb_data;
wire tile115_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile115_jtag_ucb_data;
wire tile131_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile131_jtag_ucb_data;
wire tile147_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile147_jtag_ucb_data;
wire tile163_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile163_jtag_ucb_data;
wire tile179_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile179_jtag_ucb_data;
wire tile195_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile195_jtag_ucb_data;
wire tile211_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile211_jtag_ucb_data;
wire tile227_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile227_jtag_ucb_data;
wire tile243_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile243_jtag_ucb_data;
wire tile4_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile4_jtag_ucb_data;
wire tile20_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile20_jtag_ucb_data;
wire tile36_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile36_jtag_ucb_data;
wire tile52_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile52_jtag_ucb_data;
wire tile68_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile68_jtag_ucb_data;
wire tile84_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile84_jtag_ucb_data;
wire tile100_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile100_jtag_ucb_data;
wire tile116_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile116_jtag_ucb_data;
wire tile132_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile132_jtag_ucb_data;
wire tile148_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile148_jtag_ucb_data;
wire tile164_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile164_jtag_ucb_data;
wire tile180_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile180_jtag_ucb_data;
wire tile196_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile196_jtag_ucb_data;
wire tile212_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile212_jtag_ucb_data;
wire tile228_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile228_jtag_ucb_data;
wire tile244_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile244_jtag_ucb_data;
wire tile5_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile5_jtag_ucb_data;
wire tile21_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile21_jtag_ucb_data;
wire tile37_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile37_jtag_ucb_data;
wire tile53_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile53_jtag_ucb_data;
wire tile69_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile69_jtag_ucb_data;
wire tile85_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile85_jtag_ucb_data;
wire tile101_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile101_jtag_ucb_data;
wire tile117_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile117_jtag_ucb_data;
wire tile133_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile133_jtag_ucb_data;
wire tile149_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile149_jtag_ucb_data;
wire tile165_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile165_jtag_ucb_data;
wire tile181_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile181_jtag_ucb_data;
wire tile197_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile197_jtag_ucb_data;
wire tile213_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile213_jtag_ucb_data;
wire tile229_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile229_jtag_ucb_data;
wire tile245_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile245_jtag_ucb_data;
wire tile6_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile6_jtag_ucb_data;
wire tile22_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile22_jtag_ucb_data;
wire tile38_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile38_jtag_ucb_data;
wire tile54_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile54_jtag_ucb_data;
wire tile70_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile70_jtag_ucb_data;
wire tile86_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile86_jtag_ucb_data;
wire tile102_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile102_jtag_ucb_data;
wire tile118_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile118_jtag_ucb_data;
wire tile134_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile134_jtag_ucb_data;
wire tile150_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile150_jtag_ucb_data;
wire tile166_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile166_jtag_ucb_data;
wire tile182_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile182_jtag_ucb_data;
wire tile198_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile198_jtag_ucb_data;
wire tile214_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile214_jtag_ucb_data;
wire tile230_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile230_jtag_ucb_data;
wire tile246_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile246_jtag_ucb_data;
wire tile7_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile7_jtag_ucb_data;
wire tile23_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile23_jtag_ucb_data;
wire tile39_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile39_jtag_ucb_data;
wire tile55_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile55_jtag_ucb_data;
wire tile71_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile71_jtag_ucb_data;
wire tile87_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile87_jtag_ucb_data;
wire tile103_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile103_jtag_ucb_data;
wire tile119_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile119_jtag_ucb_data;
wire tile135_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile135_jtag_ucb_data;
wire tile151_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile151_jtag_ucb_data;
wire tile167_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile167_jtag_ucb_data;
wire tile183_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile183_jtag_ucb_data;
wire tile199_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile199_jtag_ucb_data;
wire tile215_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile215_jtag_ucb_data;
wire tile231_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile231_jtag_ucb_data;
wire tile247_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile247_jtag_ucb_data;
wire tile8_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile8_jtag_ucb_data;
wire tile24_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile24_jtag_ucb_data;
wire tile40_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile40_jtag_ucb_data;
wire tile56_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile56_jtag_ucb_data;
wire tile72_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile72_jtag_ucb_data;
wire tile88_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile88_jtag_ucb_data;
wire tile104_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile104_jtag_ucb_data;
wire tile120_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile120_jtag_ucb_data;
wire tile136_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile136_jtag_ucb_data;
wire tile152_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile152_jtag_ucb_data;
wire tile168_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile168_jtag_ucb_data;
wire tile184_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile184_jtag_ucb_data;
wire tile200_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile200_jtag_ucb_data;
wire tile216_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile216_jtag_ucb_data;
wire tile232_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile232_jtag_ucb_data;
wire tile248_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile248_jtag_ucb_data;
wire tile9_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile9_jtag_ucb_data;
wire tile25_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile25_jtag_ucb_data;
wire tile41_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile41_jtag_ucb_data;
wire tile57_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile57_jtag_ucb_data;
wire tile73_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile73_jtag_ucb_data;
wire tile89_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile89_jtag_ucb_data;
wire tile105_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile105_jtag_ucb_data;
wire tile121_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile121_jtag_ucb_data;
wire tile137_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile137_jtag_ucb_data;
wire tile153_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile153_jtag_ucb_data;
wire tile169_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile169_jtag_ucb_data;
wire tile185_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile185_jtag_ucb_data;
wire tile201_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile201_jtag_ucb_data;
wire tile217_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile217_jtag_ucb_data;
wire tile233_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile233_jtag_ucb_data;
wire tile249_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile249_jtag_ucb_data;
wire tile10_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile10_jtag_ucb_data;
wire tile26_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile26_jtag_ucb_data;
wire tile42_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile42_jtag_ucb_data;
wire tile58_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile58_jtag_ucb_data;
wire tile74_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile74_jtag_ucb_data;
wire tile90_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile90_jtag_ucb_data;
wire tile106_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile106_jtag_ucb_data;
wire tile122_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile122_jtag_ucb_data;
wire tile138_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile138_jtag_ucb_data;
wire tile154_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile154_jtag_ucb_data;
wire tile170_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile170_jtag_ucb_data;
wire tile186_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile186_jtag_ucb_data;
wire tile202_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile202_jtag_ucb_data;
wire tile218_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile218_jtag_ucb_data;
wire tile234_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile234_jtag_ucb_data;
wire tile250_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile250_jtag_ucb_data;
wire tile11_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile11_jtag_ucb_data;
wire tile27_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile27_jtag_ucb_data;
wire tile43_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile43_jtag_ucb_data;
wire tile59_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile59_jtag_ucb_data;
wire tile75_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile75_jtag_ucb_data;
wire tile91_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile91_jtag_ucb_data;
wire tile107_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile107_jtag_ucb_data;
wire tile123_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile123_jtag_ucb_data;
wire tile139_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile139_jtag_ucb_data;
wire tile155_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile155_jtag_ucb_data;
wire tile171_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile171_jtag_ucb_data;
wire tile187_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile187_jtag_ucb_data;
wire tile203_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile203_jtag_ucb_data;
wire tile219_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile219_jtag_ucb_data;
wire tile235_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile235_jtag_ucb_data;
wire tile251_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile251_jtag_ucb_data;
wire tile12_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile12_jtag_ucb_data;
wire tile28_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile28_jtag_ucb_data;
wire tile44_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile44_jtag_ucb_data;
wire tile60_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile60_jtag_ucb_data;
wire tile76_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile76_jtag_ucb_data;
wire tile92_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile92_jtag_ucb_data;
wire tile108_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile108_jtag_ucb_data;
wire tile124_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile124_jtag_ucb_data;
wire tile140_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile140_jtag_ucb_data;
wire tile156_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile156_jtag_ucb_data;
wire tile172_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile172_jtag_ucb_data;
wire tile188_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile188_jtag_ucb_data;
wire tile204_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile204_jtag_ucb_data;
wire tile220_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile220_jtag_ucb_data;
wire tile236_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile236_jtag_ucb_data;
wire tile252_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile252_jtag_ucb_data;
wire tile13_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile13_jtag_ucb_data;
wire tile29_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile29_jtag_ucb_data;
wire tile45_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile45_jtag_ucb_data;
wire tile61_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile61_jtag_ucb_data;
wire tile77_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile77_jtag_ucb_data;
wire tile93_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile93_jtag_ucb_data;
wire tile109_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile109_jtag_ucb_data;
wire tile125_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile125_jtag_ucb_data;
wire tile141_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile141_jtag_ucb_data;
wire tile157_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile157_jtag_ucb_data;
wire tile173_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile173_jtag_ucb_data;
wire tile189_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile189_jtag_ucb_data;
wire tile205_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile205_jtag_ucb_data;
wire tile221_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile221_jtag_ucb_data;
wire tile237_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile237_jtag_ucb_data;
wire tile253_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile253_jtag_ucb_data;
wire tile14_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile14_jtag_ucb_data;
wire tile30_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile30_jtag_ucb_data;
wire tile46_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile46_jtag_ucb_data;
wire tile62_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile62_jtag_ucb_data;
wire tile78_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile78_jtag_ucb_data;
wire tile94_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile94_jtag_ucb_data;
wire tile110_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile110_jtag_ucb_data;
wire tile126_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile126_jtag_ucb_data;
wire tile142_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile142_jtag_ucb_data;
wire tile158_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile158_jtag_ucb_data;
wire tile174_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile174_jtag_ucb_data;
wire tile190_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile190_jtag_ucb_data;
wire tile206_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile206_jtag_ucb_data;
wire tile222_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile222_jtag_ucb_data;
wire tile238_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile238_jtag_ucb_data;
wire tile254_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile254_jtag_ucb_data;
wire tile15_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile15_jtag_ucb_data;
wire tile31_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile31_jtag_ucb_data;
wire tile47_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile47_jtag_ucb_data;
wire tile63_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile63_jtag_ucb_data;
wire tile79_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile79_jtag_ucb_data;
wire tile95_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile95_jtag_ucb_data;
wire tile111_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile111_jtag_ucb_data;
wire tile127_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile127_jtag_ucb_data;
wire tile143_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile143_jtag_ucb_data;
wire tile159_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile159_jtag_ucb_data;
wire tile175_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile175_jtag_ucb_data;
wire tile191_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile191_jtag_ucb_data;
wire tile207_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile207_jtag_ucb_data;
wire tile223_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile223_jtag_ucb_data;
wire tile239_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile239_jtag_ucb_data;
wire tile255_jtag_ucb_val;
wire [`UCB_BUS_WIDTH-1:0] tile255_jtag_ucb_data;


   // Generate tile wiring
wire [`DATA_WIDTH-1:0] tile_0_0_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_0_0_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_0_0_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_0_0_out_W_noc1_data;
wire tile_0_0_out_N_noc1_valid;
wire tile_0_0_out_S_noc1_valid;
wire tile_0_0_out_E_noc1_valid;
wire tile_0_0_out_W_noc1_valid;
wire tile_0_0_out_N_noc1_yummy;
wire tile_0_0_out_S_noc1_yummy;
wire tile_0_0_out_E_noc1_yummy;
wire tile_0_0_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_0_0_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_0_0_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_0_0_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_0_0_out_W_noc2_data;
wire tile_0_0_out_N_noc2_valid;
wire tile_0_0_out_S_noc2_valid;
wire tile_0_0_out_E_noc2_valid;
wire tile_0_0_out_W_noc2_valid;
wire tile_0_0_out_N_noc2_yummy;
wire tile_0_0_out_S_noc2_yummy;
wire tile_0_0_out_E_noc2_yummy;
wire tile_0_0_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_0_0_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_0_0_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_0_0_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_0_0_out_W_noc3_data;
wire tile_0_0_out_N_noc3_valid;
wire tile_0_0_out_S_noc3_valid;
wire tile_0_0_out_E_noc3_valid;
wire tile_0_0_out_W_noc3_valid;
wire tile_0_0_out_N_noc3_yummy;
wire tile_0_0_out_S_noc3_yummy;
wire tile_0_0_out_E_noc3_yummy;
wire tile_0_0_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_1_0_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_1_0_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_1_0_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_1_0_out_W_noc1_data;
wire tile_1_0_out_N_noc1_valid;
wire tile_1_0_out_S_noc1_valid;
wire tile_1_0_out_E_noc1_valid;
wire tile_1_0_out_W_noc1_valid;
wire tile_1_0_out_N_noc1_yummy;
wire tile_1_0_out_S_noc1_yummy;
wire tile_1_0_out_E_noc1_yummy;
wire tile_1_0_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_1_0_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_1_0_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_1_0_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_1_0_out_W_noc2_data;
wire tile_1_0_out_N_noc2_valid;
wire tile_1_0_out_S_noc2_valid;
wire tile_1_0_out_E_noc2_valid;
wire tile_1_0_out_W_noc2_valid;
wire tile_1_0_out_N_noc2_yummy;
wire tile_1_0_out_S_noc2_yummy;
wire tile_1_0_out_E_noc2_yummy;
wire tile_1_0_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_1_0_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_1_0_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_1_0_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_1_0_out_W_noc3_data;
wire tile_1_0_out_N_noc3_valid;
wire tile_1_0_out_S_noc3_valid;
wire tile_1_0_out_E_noc3_valid;
wire tile_1_0_out_W_noc3_valid;
wire tile_1_0_out_N_noc3_yummy;
wire tile_1_0_out_S_noc3_yummy;
wire tile_1_0_out_E_noc3_yummy;
wire tile_1_0_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_2_0_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_2_0_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_2_0_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_2_0_out_W_noc1_data;
wire tile_2_0_out_N_noc1_valid;
wire tile_2_0_out_S_noc1_valid;
wire tile_2_0_out_E_noc1_valid;
wire tile_2_0_out_W_noc1_valid;
wire tile_2_0_out_N_noc1_yummy;
wire tile_2_0_out_S_noc1_yummy;
wire tile_2_0_out_E_noc1_yummy;
wire tile_2_0_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_2_0_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_2_0_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_2_0_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_2_0_out_W_noc2_data;
wire tile_2_0_out_N_noc2_valid;
wire tile_2_0_out_S_noc2_valid;
wire tile_2_0_out_E_noc2_valid;
wire tile_2_0_out_W_noc2_valid;
wire tile_2_0_out_N_noc2_yummy;
wire tile_2_0_out_S_noc2_yummy;
wire tile_2_0_out_E_noc2_yummy;
wire tile_2_0_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_2_0_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_2_0_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_2_0_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_2_0_out_W_noc3_data;
wire tile_2_0_out_N_noc3_valid;
wire tile_2_0_out_S_noc3_valid;
wire tile_2_0_out_E_noc3_valid;
wire tile_2_0_out_W_noc3_valid;
wire tile_2_0_out_N_noc3_yummy;
wire tile_2_0_out_S_noc3_yummy;
wire tile_2_0_out_E_noc3_yummy;
wire tile_2_0_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_3_0_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_3_0_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_3_0_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_3_0_out_W_noc1_data;
wire tile_3_0_out_N_noc1_valid;
wire tile_3_0_out_S_noc1_valid;
wire tile_3_0_out_E_noc1_valid;
wire tile_3_0_out_W_noc1_valid;
wire tile_3_0_out_N_noc1_yummy;
wire tile_3_0_out_S_noc1_yummy;
wire tile_3_0_out_E_noc1_yummy;
wire tile_3_0_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_3_0_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_3_0_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_3_0_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_3_0_out_W_noc2_data;
wire tile_3_0_out_N_noc2_valid;
wire tile_3_0_out_S_noc2_valid;
wire tile_3_0_out_E_noc2_valid;
wire tile_3_0_out_W_noc2_valid;
wire tile_3_0_out_N_noc2_yummy;
wire tile_3_0_out_S_noc2_yummy;
wire tile_3_0_out_E_noc2_yummy;
wire tile_3_0_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_3_0_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_3_0_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_3_0_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_3_0_out_W_noc3_data;
wire tile_3_0_out_N_noc3_valid;
wire tile_3_0_out_S_noc3_valid;
wire tile_3_0_out_E_noc3_valid;
wire tile_3_0_out_W_noc3_valid;
wire tile_3_0_out_N_noc3_yummy;
wire tile_3_0_out_S_noc3_yummy;
wire tile_3_0_out_E_noc3_yummy;
wire tile_3_0_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_4_0_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_4_0_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_4_0_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_4_0_out_W_noc1_data;
wire tile_4_0_out_N_noc1_valid;
wire tile_4_0_out_S_noc1_valid;
wire tile_4_0_out_E_noc1_valid;
wire tile_4_0_out_W_noc1_valid;
wire tile_4_0_out_N_noc1_yummy;
wire tile_4_0_out_S_noc1_yummy;
wire tile_4_0_out_E_noc1_yummy;
wire tile_4_0_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_4_0_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_4_0_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_4_0_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_4_0_out_W_noc2_data;
wire tile_4_0_out_N_noc2_valid;
wire tile_4_0_out_S_noc2_valid;
wire tile_4_0_out_E_noc2_valid;
wire tile_4_0_out_W_noc2_valid;
wire tile_4_0_out_N_noc2_yummy;
wire tile_4_0_out_S_noc2_yummy;
wire tile_4_0_out_E_noc2_yummy;
wire tile_4_0_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_4_0_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_4_0_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_4_0_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_4_0_out_W_noc3_data;
wire tile_4_0_out_N_noc3_valid;
wire tile_4_0_out_S_noc3_valid;
wire tile_4_0_out_E_noc3_valid;
wire tile_4_0_out_W_noc3_valid;
wire tile_4_0_out_N_noc3_yummy;
wire tile_4_0_out_S_noc3_yummy;
wire tile_4_0_out_E_noc3_yummy;
wire tile_4_0_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_5_0_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_5_0_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_5_0_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_5_0_out_W_noc1_data;
wire tile_5_0_out_N_noc1_valid;
wire tile_5_0_out_S_noc1_valid;
wire tile_5_0_out_E_noc1_valid;
wire tile_5_0_out_W_noc1_valid;
wire tile_5_0_out_N_noc1_yummy;
wire tile_5_0_out_S_noc1_yummy;
wire tile_5_0_out_E_noc1_yummy;
wire tile_5_0_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_5_0_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_5_0_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_5_0_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_5_0_out_W_noc2_data;
wire tile_5_0_out_N_noc2_valid;
wire tile_5_0_out_S_noc2_valid;
wire tile_5_0_out_E_noc2_valid;
wire tile_5_0_out_W_noc2_valid;
wire tile_5_0_out_N_noc2_yummy;
wire tile_5_0_out_S_noc2_yummy;
wire tile_5_0_out_E_noc2_yummy;
wire tile_5_0_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_5_0_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_5_0_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_5_0_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_5_0_out_W_noc3_data;
wire tile_5_0_out_N_noc3_valid;
wire tile_5_0_out_S_noc3_valid;
wire tile_5_0_out_E_noc3_valid;
wire tile_5_0_out_W_noc3_valid;
wire tile_5_0_out_N_noc3_yummy;
wire tile_5_0_out_S_noc3_yummy;
wire tile_5_0_out_E_noc3_yummy;
wire tile_5_0_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_6_0_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_6_0_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_6_0_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_6_0_out_W_noc1_data;
wire tile_6_0_out_N_noc1_valid;
wire tile_6_0_out_S_noc1_valid;
wire tile_6_0_out_E_noc1_valid;
wire tile_6_0_out_W_noc1_valid;
wire tile_6_0_out_N_noc1_yummy;
wire tile_6_0_out_S_noc1_yummy;
wire tile_6_0_out_E_noc1_yummy;
wire tile_6_0_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_6_0_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_6_0_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_6_0_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_6_0_out_W_noc2_data;
wire tile_6_0_out_N_noc2_valid;
wire tile_6_0_out_S_noc2_valid;
wire tile_6_0_out_E_noc2_valid;
wire tile_6_0_out_W_noc2_valid;
wire tile_6_0_out_N_noc2_yummy;
wire tile_6_0_out_S_noc2_yummy;
wire tile_6_0_out_E_noc2_yummy;
wire tile_6_0_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_6_0_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_6_0_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_6_0_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_6_0_out_W_noc3_data;
wire tile_6_0_out_N_noc3_valid;
wire tile_6_0_out_S_noc3_valid;
wire tile_6_0_out_E_noc3_valid;
wire tile_6_0_out_W_noc3_valid;
wire tile_6_0_out_N_noc3_yummy;
wire tile_6_0_out_S_noc3_yummy;
wire tile_6_0_out_E_noc3_yummy;
wire tile_6_0_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_7_0_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_7_0_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_7_0_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_7_0_out_W_noc1_data;
wire tile_7_0_out_N_noc1_valid;
wire tile_7_0_out_S_noc1_valid;
wire tile_7_0_out_E_noc1_valid;
wire tile_7_0_out_W_noc1_valid;
wire tile_7_0_out_N_noc1_yummy;
wire tile_7_0_out_S_noc1_yummy;
wire tile_7_0_out_E_noc1_yummy;
wire tile_7_0_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_7_0_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_7_0_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_7_0_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_7_0_out_W_noc2_data;
wire tile_7_0_out_N_noc2_valid;
wire tile_7_0_out_S_noc2_valid;
wire tile_7_0_out_E_noc2_valid;
wire tile_7_0_out_W_noc2_valid;
wire tile_7_0_out_N_noc2_yummy;
wire tile_7_0_out_S_noc2_yummy;
wire tile_7_0_out_E_noc2_yummy;
wire tile_7_0_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_7_0_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_7_0_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_7_0_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_7_0_out_W_noc3_data;
wire tile_7_0_out_N_noc3_valid;
wire tile_7_0_out_S_noc3_valid;
wire tile_7_0_out_E_noc3_valid;
wire tile_7_0_out_W_noc3_valid;
wire tile_7_0_out_N_noc3_yummy;
wire tile_7_0_out_S_noc3_yummy;
wire tile_7_0_out_E_noc3_yummy;
wire tile_7_0_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_8_0_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_8_0_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_8_0_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_8_0_out_W_noc1_data;
wire tile_8_0_out_N_noc1_valid;
wire tile_8_0_out_S_noc1_valid;
wire tile_8_0_out_E_noc1_valid;
wire tile_8_0_out_W_noc1_valid;
wire tile_8_0_out_N_noc1_yummy;
wire tile_8_0_out_S_noc1_yummy;
wire tile_8_0_out_E_noc1_yummy;
wire tile_8_0_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_8_0_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_8_0_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_8_0_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_8_0_out_W_noc2_data;
wire tile_8_0_out_N_noc2_valid;
wire tile_8_0_out_S_noc2_valid;
wire tile_8_0_out_E_noc2_valid;
wire tile_8_0_out_W_noc2_valid;
wire tile_8_0_out_N_noc2_yummy;
wire tile_8_0_out_S_noc2_yummy;
wire tile_8_0_out_E_noc2_yummy;
wire tile_8_0_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_8_0_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_8_0_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_8_0_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_8_0_out_W_noc3_data;
wire tile_8_0_out_N_noc3_valid;
wire tile_8_0_out_S_noc3_valid;
wire tile_8_0_out_E_noc3_valid;
wire tile_8_0_out_W_noc3_valid;
wire tile_8_0_out_N_noc3_yummy;
wire tile_8_0_out_S_noc3_yummy;
wire tile_8_0_out_E_noc3_yummy;
wire tile_8_0_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_9_0_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_9_0_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_9_0_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_9_0_out_W_noc1_data;
wire tile_9_0_out_N_noc1_valid;
wire tile_9_0_out_S_noc1_valid;
wire tile_9_0_out_E_noc1_valid;
wire tile_9_0_out_W_noc1_valid;
wire tile_9_0_out_N_noc1_yummy;
wire tile_9_0_out_S_noc1_yummy;
wire tile_9_0_out_E_noc1_yummy;
wire tile_9_0_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_9_0_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_9_0_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_9_0_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_9_0_out_W_noc2_data;
wire tile_9_0_out_N_noc2_valid;
wire tile_9_0_out_S_noc2_valid;
wire tile_9_0_out_E_noc2_valid;
wire tile_9_0_out_W_noc2_valid;
wire tile_9_0_out_N_noc2_yummy;
wire tile_9_0_out_S_noc2_yummy;
wire tile_9_0_out_E_noc2_yummy;
wire tile_9_0_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_9_0_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_9_0_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_9_0_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_9_0_out_W_noc3_data;
wire tile_9_0_out_N_noc3_valid;
wire tile_9_0_out_S_noc3_valid;
wire tile_9_0_out_E_noc3_valid;
wire tile_9_0_out_W_noc3_valid;
wire tile_9_0_out_N_noc3_yummy;
wire tile_9_0_out_S_noc3_yummy;
wire tile_9_0_out_E_noc3_yummy;
wire tile_9_0_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_10_0_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_10_0_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_10_0_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_10_0_out_W_noc1_data;
wire tile_10_0_out_N_noc1_valid;
wire tile_10_0_out_S_noc1_valid;
wire tile_10_0_out_E_noc1_valid;
wire tile_10_0_out_W_noc1_valid;
wire tile_10_0_out_N_noc1_yummy;
wire tile_10_0_out_S_noc1_yummy;
wire tile_10_0_out_E_noc1_yummy;
wire tile_10_0_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_10_0_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_10_0_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_10_0_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_10_0_out_W_noc2_data;
wire tile_10_0_out_N_noc2_valid;
wire tile_10_0_out_S_noc2_valid;
wire tile_10_0_out_E_noc2_valid;
wire tile_10_0_out_W_noc2_valid;
wire tile_10_0_out_N_noc2_yummy;
wire tile_10_0_out_S_noc2_yummy;
wire tile_10_0_out_E_noc2_yummy;
wire tile_10_0_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_10_0_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_10_0_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_10_0_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_10_0_out_W_noc3_data;
wire tile_10_0_out_N_noc3_valid;
wire tile_10_0_out_S_noc3_valid;
wire tile_10_0_out_E_noc3_valid;
wire tile_10_0_out_W_noc3_valid;
wire tile_10_0_out_N_noc3_yummy;
wire tile_10_0_out_S_noc3_yummy;
wire tile_10_0_out_E_noc3_yummy;
wire tile_10_0_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_11_0_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_11_0_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_11_0_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_11_0_out_W_noc1_data;
wire tile_11_0_out_N_noc1_valid;
wire tile_11_0_out_S_noc1_valid;
wire tile_11_0_out_E_noc1_valid;
wire tile_11_0_out_W_noc1_valid;
wire tile_11_0_out_N_noc1_yummy;
wire tile_11_0_out_S_noc1_yummy;
wire tile_11_0_out_E_noc1_yummy;
wire tile_11_0_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_11_0_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_11_0_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_11_0_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_11_0_out_W_noc2_data;
wire tile_11_0_out_N_noc2_valid;
wire tile_11_0_out_S_noc2_valid;
wire tile_11_0_out_E_noc2_valid;
wire tile_11_0_out_W_noc2_valid;
wire tile_11_0_out_N_noc2_yummy;
wire tile_11_0_out_S_noc2_yummy;
wire tile_11_0_out_E_noc2_yummy;
wire tile_11_0_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_11_0_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_11_0_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_11_0_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_11_0_out_W_noc3_data;
wire tile_11_0_out_N_noc3_valid;
wire tile_11_0_out_S_noc3_valid;
wire tile_11_0_out_E_noc3_valid;
wire tile_11_0_out_W_noc3_valid;
wire tile_11_0_out_N_noc3_yummy;
wire tile_11_0_out_S_noc3_yummy;
wire tile_11_0_out_E_noc3_yummy;
wire tile_11_0_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_12_0_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_12_0_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_12_0_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_12_0_out_W_noc1_data;
wire tile_12_0_out_N_noc1_valid;
wire tile_12_0_out_S_noc1_valid;
wire tile_12_0_out_E_noc1_valid;
wire tile_12_0_out_W_noc1_valid;
wire tile_12_0_out_N_noc1_yummy;
wire tile_12_0_out_S_noc1_yummy;
wire tile_12_0_out_E_noc1_yummy;
wire tile_12_0_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_12_0_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_12_0_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_12_0_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_12_0_out_W_noc2_data;
wire tile_12_0_out_N_noc2_valid;
wire tile_12_0_out_S_noc2_valid;
wire tile_12_0_out_E_noc2_valid;
wire tile_12_0_out_W_noc2_valid;
wire tile_12_0_out_N_noc2_yummy;
wire tile_12_0_out_S_noc2_yummy;
wire tile_12_0_out_E_noc2_yummy;
wire tile_12_0_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_12_0_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_12_0_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_12_0_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_12_0_out_W_noc3_data;
wire tile_12_0_out_N_noc3_valid;
wire tile_12_0_out_S_noc3_valid;
wire tile_12_0_out_E_noc3_valid;
wire tile_12_0_out_W_noc3_valid;
wire tile_12_0_out_N_noc3_yummy;
wire tile_12_0_out_S_noc3_yummy;
wire tile_12_0_out_E_noc3_yummy;
wire tile_12_0_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_13_0_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_13_0_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_13_0_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_13_0_out_W_noc1_data;
wire tile_13_0_out_N_noc1_valid;
wire tile_13_0_out_S_noc1_valid;
wire tile_13_0_out_E_noc1_valid;
wire tile_13_0_out_W_noc1_valid;
wire tile_13_0_out_N_noc1_yummy;
wire tile_13_0_out_S_noc1_yummy;
wire tile_13_0_out_E_noc1_yummy;
wire tile_13_0_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_13_0_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_13_0_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_13_0_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_13_0_out_W_noc2_data;
wire tile_13_0_out_N_noc2_valid;
wire tile_13_0_out_S_noc2_valid;
wire tile_13_0_out_E_noc2_valid;
wire tile_13_0_out_W_noc2_valid;
wire tile_13_0_out_N_noc2_yummy;
wire tile_13_0_out_S_noc2_yummy;
wire tile_13_0_out_E_noc2_yummy;
wire tile_13_0_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_13_0_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_13_0_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_13_0_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_13_0_out_W_noc3_data;
wire tile_13_0_out_N_noc3_valid;
wire tile_13_0_out_S_noc3_valid;
wire tile_13_0_out_E_noc3_valid;
wire tile_13_0_out_W_noc3_valid;
wire tile_13_0_out_N_noc3_yummy;
wire tile_13_0_out_S_noc3_yummy;
wire tile_13_0_out_E_noc3_yummy;
wire tile_13_0_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_14_0_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_14_0_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_14_0_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_14_0_out_W_noc1_data;
wire tile_14_0_out_N_noc1_valid;
wire tile_14_0_out_S_noc1_valid;
wire tile_14_0_out_E_noc1_valid;
wire tile_14_0_out_W_noc1_valid;
wire tile_14_0_out_N_noc1_yummy;
wire tile_14_0_out_S_noc1_yummy;
wire tile_14_0_out_E_noc1_yummy;
wire tile_14_0_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_14_0_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_14_0_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_14_0_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_14_0_out_W_noc2_data;
wire tile_14_0_out_N_noc2_valid;
wire tile_14_0_out_S_noc2_valid;
wire tile_14_0_out_E_noc2_valid;
wire tile_14_0_out_W_noc2_valid;
wire tile_14_0_out_N_noc2_yummy;
wire tile_14_0_out_S_noc2_yummy;
wire tile_14_0_out_E_noc2_yummy;
wire tile_14_0_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_14_0_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_14_0_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_14_0_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_14_0_out_W_noc3_data;
wire tile_14_0_out_N_noc3_valid;
wire tile_14_0_out_S_noc3_valid;
wire tile_14_0_out_E_noc3_valid;
wire tile_14_0_out_W_noc3_valid;
wire tile_14_0_out_N_noc3_yummy;
wire tile_14_0_out_S_noc3_yummy;
wire tile_14_0_out_E_noc3_yummy;
wire tile_14_0_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_15_0_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_15_0_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_15_0_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_15_0_out_W_noc1_data;
wire tile_15_0_out_N_noc1_valid;
wire tile_15_0_out_S_noc1_valid;
wire tile_15_0_out_E_noc1_valid;
wire tile_15_0_out_W_noc1_valid;
wire tile_15_0_out_N_noc1_yummy;
wire tile_15_0_out_S_noc1_yummy;
wire tile_15_0_out_E_noc1_yummy;
wire tile_15_0_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_15_0_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_15_0_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_15_0_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_15_0_out_W_noc2_data;
wire tile_15_0_out_N_noc2_valid;
wire tile_15_0_out_S_noc2_valid;
wire tile_15_0_out_E_noc2_valid;
wire tile_15_0_out_W_noc2_valid;
wire tile_15_0_out_N_noc2_yummy;
wire tile_15_0_out_S_noc2_yummy;
wire tile_15_0_out_E_noc2_yummy;
wire tile_15_0_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_15_0_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_15_0_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_15_0_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_15_0_out_W_noc3_data;
wire tile_15_0_out_N_noc3_valid;
wire tile_15_0_out_S_noc3_valid;
wire tile_15_0_out_E_noc3_valid;
wire tile_15_0_out_W_noc3_valid;
wire tile_15_0_out_N_noc3_yummy;
wire tile_15_0_out_S_noc3_yummy;
wire tile_15_0_out_E_noc3_yummy;
wire tile_15_0_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_0_1_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_0_1_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_0_1_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_0_1_out_W_noc1_data;
wire tile_0_1_out_N_noc1_valid;
wire tile_0_1_out_S_noc1_valid;
wire tile_0_1_out_E_noc1_valid;
wire tile_0_1_out_W_noc1_valid;
wire tile_0_1_out_N_noc1_yummy;
wire tile_0_1_out_S_noc1_yummy;
wire tile_0_1_out_E_noc1_yummy;
wire tile_0_1_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_0_1_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_0_1_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_0_1_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_0_1_out_W_noc2_data;
wire tile_0_1_out_N_noc2_valid;
wire tile_0_1_out_S_noc2_valid;
wire tile_0_1_out_E_noc2_valid;
wire tile_0_1_out_W_noc2_valid;
wire tile_0_1_out_N_noc2_yummy;
wire tile_0_1_out_S_noc2_yummy;
wire tile_0_1_out_E_noc2_yummy;
wire tile_0_1_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_0_1_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_0_1_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_0_1_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_0_1_out_W_noc3_data;
wire tile_0_1_out_N_noc3_valid;
wire tile_0_1_out_S_noc3_valid;
wire tile_0_1_out_E_noc3_valid;
wire tile_0_1_out_W_noc3_valid;
wire tile_0_1_out_N_noc3_yummy;
wire tile_0_1_out_S_noc3_yummy;
wire tile_0_1_out_E_noc3_yummy;
wire tile_0_1_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_1_1_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_1_1_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_1_1_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_1_1_out_W_noc1_data;
wire tile_1_1_out_N_noc1_valid;
wire tile_1_1_out_S_noc1_valid;
wire tile_1_1_out_E_noc1_valid;
wire tile_1_1_out_W_noc1_valid;
wire tile_1_1_out_N_noc1_yummy;
wire tile_1_1_out_S_noc1_yummy;
wire tile_1_1_out_E_noc1_yummy;
wire tile_1_1_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_1_1_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_1_1_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_1_1_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_1_1_out_W_noc2_data;
wire tile_1_1_out_N_noc2_valid;
wire tile_1_1_out_S_noc2_valid;
wire tile_1_1_out_E_noc2_valid;
wire tile_1_1_out_W_noc2_valid;
wire tile_1_1_out_N_noc2_yummy;
wire tile_1_1_out_S_noc2_yummy;
wire tile_1_1_out_E_noc2_yummy;
wire tile_1_1_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_1_1_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_1_1_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_1_1_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_1_1_out_W_noc3_data;
wire tile_1_1_out_N_noc3_valid;
wire tile_1_1_out_S_noc3_valid;
wire tile_1_1_out_E_noc3_valid;
wire tile_1_1_out_W_noc3_valid;
wire tile_1_1_out_N_noc3_yummy;
wire tile_1_1_out_S_noc3_yummy;
wire tile_1_1_out_E_noc3_yummy;
wire tile_1_1_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_2_1_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_2_1_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_2_1_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_2_1_out_W_noc1_data;
wire tile_2_1_out_N_noc1_valid;
wire tile_2_1_out_S_noc1_valid;
wire tile_2_1_out_E_noc1_valid;
wire tile_2_1_out_W_noc1_valid;
wire tile_2_1_out_N_noc1_yummy;
wire tile_2_1_out_S_noc1_yummy;
wire tile_2_1_out_E_noc1_yummy;
wire tile_2_1_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_2_1_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_2_1_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_2_1_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_2_1_out_W_noc2_data;
wire tile_2_1_out_N_noc2_valid;
wire tile_2_1_out_S_noc2_valid;
wire tile_2_1_out_E_noc2_valid;
wire tile_2_1_out_W_noc2_valid;
wire tile_2_1_out_N_noc2_yummy;
wire tile_2_1_out_S_noc2_yummy;
wire tile_2_1_out_E_noc2_yummy;
wire tile_2_1_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_2_1_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_2_1_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_2_1_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_2_1_out_W_noc3_data;
wire tile_2_1_out_N_noc3_valid;
wire tile_2_1_out_S_noc3_valid;
wire tile_2_1_out_E_noc3_valid;
wire tile_2_1_out_W_noc3_valid;
wire tile_2_1_out_N_noc3_yummy;
wire tile_2_1_out_S_noc3_yummy;
wire tile_2_1_out_E_noc3_yummy;
wire tile_2_1_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_3_1_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_3_1_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_3_1_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_3_1_out_W_noc1_data;
wire tile_3_1_out_N_noc1_valid;
wire tile_3_1_out_S_noc1_valid;
wire tile_3_1_out_E_noc1_valid;
wire tile_3_1_out_W_noc1_valid;
wire tile_3_1_out_N_noc1_yummy;
wire tile_3_1_out_S_noc1_yummy;
wire tile_3_1_out_E_noc1_yummy;
wire tile_3_1_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_3_1_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_3_1_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_3_1_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_3_1_out_W_noc2_data;
wire tile_3_1_out_N_noc2_valid;
wire tile_3_1_out_S_noc2_valid;
wire tile_3_1_out_E_noc2_valid;
wire tile_3_1_out_W_noc2_valid;
wire tile_3_1_out_N_noc2_yummy;
wire tile_3_1_out_S_noc2_yummy;
wire tile_3_1_out_E_noc2_yummy;
wire tile_3_1_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_3_1_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_3_1_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_3_1_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_3_1_out_W_noc3_data;
wire tile_3_1_out_N_noc3_valid;
wire tile_3_1_out_S_noc3_valid;
wire tile_3_1_out_E_noc3_valid;
wire tile_3_1_out_W_noc3_valid;
wire tile_3_1_out_N_noc3_yummy;
wire tile_3_1_out_S_noc3_yummy;
wire tile_3_1_out_E_noc3_yummy;
wire tile_3_1_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_4_1_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_4_1_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_4_1_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_4_1_out_W_noc1_data;
wire tile_4_1_out_N_noc1_valid;
wire tile_4_1_out_S_noc1_valid;
wire tile_4_1_out_E_noc1_valid;
wire tile_4_1_out_W_noc1_valid;
wire tile_4_1_out_N_noc1_yummy;
wire tile_4_1_out_S_noc1_yummy;
wire tile_4_1_out_E_noc1_yummy;
wire tile_4_1_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_4_1_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_4_1_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_4_1_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_4_1_out_W_noc2_data;
wire tile_4_1_out_N_noc2_valid;
wire tile_4_1_out_S_noc2_valid;
wire tile_4_1_out_E_noc2_valid;
wire tile_4_1_out_W_noc2_valid;
wire tile_4_1_out_N_noc2_yummy;
wire tile_4_1_out_S_noc2_yummy;
wire tile_4_1_out_E_noc2_yummy;
wire tile_4_1_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_4_1_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_4_1_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_4_1_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_4_1_out_W_noc3_data;
wire tile_4_1_out_N_noc3_valid;
wire tile_4_1_out_S_noc3_valid;
wire tile_4_1_out_E_noc3_valid;
wire tile_4_1_out_W_noc3_valid;
wire tile_4_1_out_N_noc3_yummy;
wire tile_4_1_out_S_noc3_yummy;
wire tile_4_1_out_E_noc3_yummy;
wire tile_4_1_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_5_1_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_5_1_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_5_1_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_5_1_out_W_noc1_data;
wire tile_5_1_out_N_noc1_valid;
wire tile_5_1_out_S_noc1_valid;
wire tile_5_1_out_E_noc1_valid;
wire tile_5_1_out_W_noc1_valid;
wire tile_5_1_out_N_noc1_yummy;
wire tile_5_1_out_S_noc1_yummy;
wire tile_5_1_out_E_noc1_yummy;
wire tile_5_1_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_5_1_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_5_1_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_5_1_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_5_1_out_W_noc2_data;
wire tile_5_1_out_N_noc2_valid;
wire tile_5_1_out_S_noc2_valid;
wire tile_5_1_out_E_noc2_valid;
wire tile_5_1_out_W_noc2_valid;
wire tile_5_1_out_N_noc2_yummy;
wire tile_5_1_out_S_noc2_yummy;
wire tile_5_1_out_E_noc2_yummy;
wire tile_5_1_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_5_1_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_5_1_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_5_1_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_5_1_out_W_noc3_data;
wire tile_5_1_out_N_noc3_valid;
wire tile_5_1_out_S_noc3_valid;
wire tile_5_1_out_E_noc3_valid;
wire tile_5_1_out_W_noc3_valid;
wire tile_5_1_out_N_noc3_yummy;
wire tile_5_1_out_S_noc3_yummy;
wire tile_5_1_out_E_noc3_yummy;
wire tile_5_1_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_6_1_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_6_1_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_6_1_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_6_1_out_W_noc1_data;
wire tile_6_1_out_N_noc1_valid;
wire tile_6_1_out_S_noc1_valid;
wire tile_6_1_out_E_noc1_valid;
wire tile_6_1_out_W_noc1_valid;
wire tile_6_1_out_N_noc1_yummy;
wire tile_6_1_out_S_noc1_yummy;
wire tile_6_1_out_E_noc1_yummy;
wire tile_6_1_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_6_1_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_6_1_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_6_1_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_6_1_out_W_noc2_data;
wire tile_6_1_out_N_noc2_valid;
wire tile_6_1_out_S_noc2_valid;
wire tile_6_1_out_E_noc2_valid;
wire tile_6_1_out_W_noc2_valid;
wire tile_6_1_out_N_noc2_yummy;
wire tile_6_1_out_S_noc2_yummy;
wire tile_6_1_out_E_noc2_yummy;
wire tile_6_1_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_6_1_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_6_1_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_6_1_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_6_1_out_W_noc3_data;
wire tile_6_1_out_N_noc3_valid;
wire tile_6_1_out_S_noc3_valid;
wire tile_6_1_out_E_noc3_valid;
wire tile_6_1_out_W_noc3_valid;
wire tile_6_1_out_N_noc3_yummy;
wire tile_6_1_out_S_noc3_yummy;
wire tile_6_1_out_E_noc3_yummy;
wire tile_6_1_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_7_1_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_7_1_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_7_1_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_7_1_out_W_noc1_data;
wire tile_7_1_out_N_noc1_valid;
wire tile_7_1_out_S_noc1_valid;
wire tile_7_1_out_E_noc1_valid;
wire tile_7_1_out_W_noc1_valid;
wire tile_7_1_out_N_noc1_yummy;
wire tile_7_1_out_S_noc1_yummy;
wire tile_7_1_out_E_noc1_yummy;
wire tile_7_1_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_7_1_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_7_1_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_7_1_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_7_1_out_W_noc2_data;
wire tile_7_1_out_N_noc2_valid;
wire tile_7_1_out_S_noc2_valid;
wire tile_7_1_out_E_noc2_valid;
wire tile_7_1_out_W_noc2_valid;
wire tile_7_1_out_N_noc2_yummy;
wire tile_7_1_out_S_noc2_yummy;
wire tile_7_1_out_E_noc2_yummy;
wire tile_7_1_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_7_1_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_7_1_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_7_1_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_7_1_out_W_noc3_data;
wire tile_7_1_out_N_noc3_valid;
wire tile_7_1_out_S_noc3_valid;
wire tile_7_1_out_E_noc3_valid;
wire tile_7_1_out_W_noc3_valid;
wire tile_7_1_out_N_noc3_yummy;
wire tile_7_1_out_S_noc3_yummy;
wire tile_7_1_out_E_noc3_yummy;
wire tile_7_1_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_8_1_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_8_1_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_8_1_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_8_1_out_W_noc1_data;
wire tile_8_1_out_N_noc1_valid;
wire tile_8_1_out_S_noc1_valid;
wire tile_8_1_out_E_noc1_valid;
wire tile_8_1_out_W_noc1_valid;
wire tile_8_1_out_N_noc1_yummy;
wire tile_8_1_out_S_noc1_yummy;
wire tile_8_1_out_E_noc1_yummy;
wire tile_8_1_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_8_1_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_8_1_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_8_1_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_8_1_out_W_noc2_data;
wire tile_8_1_out_N_noc2_valid;
wire tile_8_1_out_S_noc2_valid;
wire tile_8_1_out_E_noc2_valid;
wire tile_8_1_out_W_noc2_valid;
wire tile_8_1_out_N_noc2_yummy;
wire tile_8_1_out_S_noc2_yummy;
wire tile_8_1_out_E_noc2_yummy;
wire tile_8_1_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_8_1_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_8_1_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_8_1_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_8_1_out_W_noc3_data;
wire tile_8_1_out_N_noc3_valid;
wire tile_8_1_out_S_noc3_valid;
wire tile_8_1_out_E_noc3_valid;
wire tile_8_1_out_W_noc3_valid;
wire tile_8_1_out_N_noc3_yummy;
wire tile_8_1_out_S_noc3_yummy;
wire tile_8_1_out_E_noc3_yummy;
wire tile_8_1_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_9_1_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_9_1_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_9_1_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_9_1_out_W_noc1_data;
wire tile_9_1_out_N_noc1_valid;
wire tile_9_1_out_S_noc1_valid;
wire tile_9_1_out_E_noc1_valid;
wire tile_9_1_out_W_noc1_valid;
wire tile_9_1_out_N_noc1_yummy;
wire tile_9_1_out_S_noc1_yummy;
wire tile_9_1_out_E_noc1_yummy;
wire tile_9_1_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_9_1_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_9_1_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_9_1_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_9_1_out_W_noc2_data;
wire tile_9_1_out_N_noc2_valid;
wire tile_9_1_out_S_noc2_valid;
wire tile_9_1_out_E_noc2_valid;
wire tile_9_1_out_W_noc2_valid;
wire tile_9_1_out_N_noc2_yummy;
wire tile_9_1_out_S_noc2_yummy;
wire tile_9_1_out_E_noc2_yummy;
wire tile_9_1_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_9_1_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_9_1_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_9_1_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_9_1_out_W_noc3_data;
wire tile_9_1_out_N_noc3_valid;
wire tile_9_1_out_S_noc3_valid;
wire tile_9_1_out_E_noc3_valid;
wire tile_9_1_out_W_noc3_valid;
wire tile_9_1_out_N_noc3_yummy;
wire tile_9_1_out_S_noc3_yummy;
wire tile_9_1_out_E_noc3_yummy;
wire tile_9_1_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_10_1_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_10_1_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_10_1_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_10_1_out_W_noc1_data;
wire tile_10_1_out_N_noc1_valid;
wire tile_10_1_out_S_noc1_valid;
wire tile_10_1_out_E_noc1_valid;
wire tile_10_1_out_W_noc1_valid;
wire tile_10_1_out_N_noc1_yummy;
wire tile_10_1_out_S_noc1_yummy;
wire tile_10_1_out_E_noc1_yummy;
wire tile_10_1_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_10_1_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_10_1_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_10_1_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_10_1_out_W_noc2_data;
wire tile_10_1_out_N_noc2_valid;
wire tile_10_1_out_S_noc2_valid;
wire tile_10_1_out_E_noc2_valid;
wire tile_10_1_out_W_noc2_valid;
wire tile_10_1_out_N_noc2_yummy;
wire tile_10_1_out_S_noc2_yummy;
wire tile_10_1_out_E_noc2_yummy;
wire tile_10_1_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_10_1_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_10_1_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_10_1_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_10_1_out_W_noc3_data;
wire tile_10_1_out_N_noc3_valid;
wire tile_10_1_out_S_noc3_valid;
wire tile_10_1_out_E_noc3_valid;
wire tile_10_1_out_W_noc3_valid;
wire tile_10_1_out_N_noc3_yummy;
wire tile_10_1_out_S_noc3_yummy;
wire tile_10_1_out_E_noc3_yummy;
wire tile_10_1_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_11_1_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_11_1_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_11_1_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_11_1_out_W_noc1_data;
wire tile_11_1_out_N_noc1_valid;
wire tile_11_1_out_S_noc1_valid;
wire tile_11_1_out_E_noc1_valid;
wire tile_11_1_out_W_noc1_valid;
wire tile_11_1_out_N_noc1_yummy;
wire tile_11_1_out_S_noc1_yummy;
wire tile_11_1_out_E_noc1_yummy;
wire tile_11_1_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_11_1_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_11_1_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_11_1_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_11_1_out_W_noc2_data;
wire tile_11_1_out_N_noc2_valid;
wire tile_11_1_out_S_noc2_valid;
wire tile_11_1_out_E_noc2_valid;
wire tile_11_1_out_W_noc2_valid;
wire tile_11_1_out_N_noc2_yummy;
wire tile_11_1_out_S_noc2_yummy;
wire tile_11_1_out_E_noc2_yummy;
wire tile_11_1_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_11_1_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_11_1_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_11_1_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_11_1_out_W_noc3_data;
wire tile_11_1_out_N_noc3_valid;
wire tile_11_1_out_S_noc3_valid;
wire tile_11_1_out_E_noc3_valid;
wire tile_11_1_out_W_noc3_valid;
wire tile_11_1_out_N_noc3_yummy;
wire tile_11_1_out_S_noc3_yummy;
wire tile_11_1_out_E_noc3_yummy;
wire tile_11_1_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_12_1_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_12_1_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_12_1_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_12_1_out_W_noc1_data;
wire tile_12_1_out_N_noc1_valid;
wire tile_12_1_out_S_noc1_valid;
wire tile_12_1_out_E_noc1_valid;
wire tile_12_1_out_W_noc1_valid;
wire tile_12_1_out_N_noc1_yummy;
wire tile_12_1_out_S_noc1_yummy;
wire tile_12_1_out_E_noc1_yummy;
wire tile_12_1_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_12_1_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_12_1_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_12_1_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_12_1_out_W_noc2_data;
wire tile_12_1_out_N_noc2_valid;
wire tile_12_1_out_S_noc2_valid;
wire tile_12_1_out_E_noc2_valid;
wire tile_12_1_out_W_noc2_valid;
wire tile_12_1_out_N_noc2_yummy;
wire tile_12_1_out_S_noc2_yummy;
wire tile_12_1_out_E_noc2_yummy;
wire tile_12_1_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_12_1_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_12_1_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_12_1_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_12_1_out_W_noc3_data;
wire tile_12_1_out_N_noc3_valid;
wire tile_12_1_out_S_noc3_valid;
wire tile_12_1_out_E_noc3_valid;
wire tile_12_1_out_W_noc3_valid;
wire tile_12_1_out_N_noc3_yummy;
wire tile_12_1_out_S_noc3_yummy;
wire tile_12_1_out_E_noc3_yummy;
wire tile_12_1_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_13_1_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_13_1_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_13_1_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_13_1_out_W_noc1_data;
wire tile_13_1_out_N_noc1_valid;
wire tile_13_1_out_S_noc1_valid;
wire tile_13_1_out_E_noc1_valid;
wire tile_13_1_out_W_noc1_valid;
wire tile_13_1_out_N_noc1_yummy;
wire tile_13_1_out_S_noc1_yummy;
wire tile_13_1_out_E_noc1_yummy;
wire tile_13_1_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_13_1_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_13_1_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_13_1_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_13_1_out_W_noc2_data;
wire tile_13_1_out_N_noc2_valid;
wire tile_13_1_out_S_noc2_valid;
wire tile_13_1_out_E_noc2_valid;
wire tile_13_1_out_W_noc2_valid;
wire tile_13_1_out_N_noc2_yummy;
wire tile_13_1_out_S_noc2_yummy;
wire tile_13_1_out_E_noc2_yummy;
wire tile_13_1_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_13_1_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_13_1_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_13_1_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_13_1_out_W_noc3_data;
wire tile_13_1_out_N_noc3_valid;
wire tile_13_1_out_S_noc3_valid;
wire tile_13_1_out_E_noc3_valid;
wire tile_13_1_out_W_noc3_valid;
wire tile_13_1_out_N_noc3_yummy;
wire tile_13_1_out_S_noc3_yummy;
wire tile_13_1_out_E_noc3_yummy;
wire tile_13_1_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_14_1_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_14_1_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_14_1_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_14_1_out_W_noc1_data;
wire tile_14_1_out_N_noc1_valid;
wire tile_14_1_out_S_noc1_valid;
wire tile_14_1_out_E_noc1_valid;
wire tile_14_1_out_W_noc1_valid;
wire tile_14_1_out_N_noc1_yummy;
wire tile_14_1_out_S_noc1_yummy;
wire tile_14_1_out_E_noc1_yummy;
wire tile_14_1_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_14_1_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_14_1_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_14_1_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_14_1_out_W_noc2_data;
wire tile_14_1_out_N_noc2_valid;
wire tile_14_1_out_S_noc2_valid;
wire tile_14_1_out_E_noc2_valid;
wire tile_14_1_out_W_noc2_valid;
wire tile_14_1_out_N_noc2_yummy;
wire tile_14_1_out_S_noc2_yummy;
wire tile_14_1_out_E_noc2_yummy;
wire tile_14_1_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_14_1_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_14_1_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_14_1_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_14_1_out_W_noc3_data;
wire tile_14_1_out_N_noc3_valid;
wire tile_14_1_out_S_noc3_valid;
wire tile_14_1_out_E_noc3_valid;
wire tile_14_1_out_W_noc3_valid;
wire tile_14_1_out_N_noc3_yummy;
wire tile_14_1_out_S_noc3_yummy;
wire tile_14_1_out_E_noc3_yummy;
wire tile_14_1_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_15_1_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_15_1_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_15_1_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_15_1_out_W_noc1_data;
wire tile_15_1_out_N_noc1_valid;
wire tile_15_1_out_S_noc1_valid;
wire tile_15_1_out_E_noc1_valid;
wire tile_15_1_out_W_noc1_valid;
wire tile_15_1_out_N_noc1_yummy;
wire tile_15_1_out_S_noc1_yummy;
wire tile_15_1_out_E_noc1_yummy;
wire tile_15_1_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_15_1_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_15_1_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_15_1_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_15_1_out_W_noc2_data;
wire tile_15_1_out_N_noc2_valid;
wire tile_15_1_out_S_noc2_valid;
wire tile_15_1_out_E_noc2_valid;
wire tile_15_1_out_W_noc2_valid;
wire tile_15_1_out_N_noc2_yummy;
wire tile_15_1_out_S_noc2_yummy;
wire tile_15_1_out_E_noc2_yummy;
wire tile_15_1_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_15_1_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_15_1_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_15_1_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_15_1_out_W_noc3_data;
wire tile_15_1_out_N_noc3_valid;
wire tile_15_1_out_S_noc3_valid;
wire tile_15_1_out_E_noc3_valid;
wire tile_15_1_out_W_noc3_valid;
wire tile_15_1_out_N_noc3_yummy;
wire tile_15_1_out_S_noc3_yummy;
wire tile_15_1_out_E_noc3_yummy;
wire tile_15_1_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_0_2_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_0_2_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_0_2_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_0_2_out_W_noc1_data;
wire tile_0_2_out_N_noc1_valid;
wire tile_0_2_out_S_noc1_valid;
wire tile_0_2_out_E_noc1_valid;
wire tile_0_2_out_W_noc1_valid;
wire tile_0_2_out_N_noc1_yummy;
wire tile_0_2_out_S_noc1_yummy;
wire tile_0_2_out_E_noc1_yummy;
wire tile_0_2_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_0_2_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_0_2_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_0_2_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_0_2_out_W_noc2_data;
wire tile_0_2_out_N_noc2_valid;
wire tile_0_2_out_S_noc2_valid;
wire tile_0_2_out_E_noc2_valid;
wire tile_0_2_out_W_noc2_valid;
wire tile_0_2_out_N_noc2_yummy;
wire tile_0_2_out_S_noc2_yummy;
wire tile_0_2_out_E_noc2_yummy;
wire tile_0_2_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_0_2_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_0_2_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_0_2_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_0_2_out_W_noc3_data;
wire tile_0_2_out_N_noc3_valid;
wire tile_0_2_out_S_noc3_valid;
wire tile_0_2_out_E_noc3_valid;
wire tile_0_2_out_W_noc3_valid;
wire tile_0_2_out_N_noc3_yummy;
wire tile_0_2_out_S_noc3_yummy;
wire tile_0_2_out_E_noc3_yummy;
wire tile_0_2_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_1_2_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_1_2_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_1_2_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_1_2_out_W_noc1_data;
wire tile_1_2_out_N_noc1_valid;
wire tile_1_2_out_S_noc1_valid;
wire tile_1_2_out_E_noc1_valid;
wire tile_1_2_out_W_noc1_valid;
wire tile_1_2_out_N_noc1_yummy;
wire tile_1_2_out_S_noc1_yummy;
wire tile_1_2_out_E_noc1_yummy;
wire tile_1_2_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_1_2_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_1_2_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_1_2_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_1_2_out_W_noc2_data;
wire tile_1_2_out_N_noc2_valid;
wire tile_1_2_out_S_noc2_valid;
wire tile_1_2_out_E_noc2_valid;
wire tile_1_2_out_W_noc2_valid;
wire tile_1_2_out_N_noc2_yummy;
wire tile_1_2_out_S_noc2_yummy;
wire tile_1_2_out_E_noc2_yummy;
wire tile_1_2_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_1_2_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_1_2_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_1_2_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_1_2_out_W_noc3_data;
wire tile_1_2_out_N_noc3_valid;
wire tile_1_2_out_S_noc3_valid;
wire tile_1_2_out_E_noc3_valid;
wire tile_1_2_out_W_noc3_valid;
wire tile_1_2_out_N_noc3_yummy;
wire tile_1_2_out_S_noc3_yummy;
wire tile_1_2_out_E_noc3_yummy;
wire tile_1_2_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_2_2_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_2_2_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_2_2_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_2_2_out_W_noc1_data;
wire tile_2_2_out_N_noc1_valid;
wire tile_2_2_out_S_noc1_valid;
wire tile_2_2_out_E_noc1_valid;
wire tile_2_2_out_W_noc1_valid;
wire tile_2_2_out_N_noc1_yummy;
wire tile_2_2_out_S_noc1_yummy;
wire tile_2_2_out_E_noc1_yummy;
wire tile_2_2_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_2_2_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_2_2_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_2_2_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_2_2_out_W_noc2_data;
wire tile_2_2_out_N_noc2_valid;
wire tile_2_2_out_S_noc2_valid;
wire tile_2_2_out_E_noc2_valid;
wire tile_2_2_out_W_noc2_valid;
wire tile_2_2_out_N_noc2_yummy;
wire tile_2_2_out_S_noc2_yummy;
wire tile_2_2_out_E_noc2_yummy;
wire tile_2_2_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_2_2_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_2_2_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_2_2_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_2_2_out_W_noc3_data;
wire tile_2_2_out_N_noc3_valid;
wire tile_2_2_out_S_noc3_valid;
wire tile_2_2_out_E_noc3_valid;
wire tile_2_2_out_W_noc3_valid;
wire tile_2_2_out_N_noc3_yummy;
wire tile_2_2_out_S_noc3_yummy;
wire tile_2_2_out_E_noc3_yummy;
wire tile_2_2_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_3_2_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_3_2_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_3_2_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_3_2_out_W_noc1_data;
wire tile_3_2_out_N_noc1_valid;
wire tile_3_2_out_S_noc1_valid;
wire tile_3_2_out_E_noc1_valid;
wire tile_3_2_out_W_noc1_valid;
wire tile_3_2_out_N_noc1_yummy;
wire tile_3_2_out_S_noc1_yummy;
wire tile_3_2_out_E_noc1_yummy;
wire tile_3_2_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_3_2_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_3_2_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_3_2_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_3_2_out_W_noc2_data;
wire tile_3_2_out_N_noc2_valid;
wire tile_3_2_out_S_noc2_valid;
wire tile_3_2_out_E_noc2_valid;
wire tile_3_2_out_W_noc2_valid;
wire tile_3_2_out_N_noc2_yummy;
wire tile_3_2_out_S_noc2_yummy;
wire tile_3_2_out_E_noc2_yummy;
wire tile_3_2_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_3_2_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_3_2_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_3_2_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_3_2_out_W_noc3_data;
wire tile_3_2_out_N_noc3_valid;
wire tile_3_2_out_S_noc3_valid;
wire tile_3_2_out_E_noc3_valid;
wire tile_3_2_out_W_noc3_valid;
wire tile_3_2_out_N_noc3_yummy;
wire tile_3_2_out_S_noc3_yummy;
wire tile_3_2_out_E_noc3_yummy;
wire tile_3_2_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_4_2_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_4_2_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_4_2_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_4_2_out_W_noc1_data;
wire tile_4_2_out_N_noc1_valid;
wire tile_4_2_out_S_noc1_valid;
wire tile_4_2_out_E_noc1_valid;
wire tile_4_2_out_W_noc1_valid;
wire tile_4_2_out_N_noc1_yummy;
wire tile_4_2_out_S_noc1_yummy;
wire tile_4_2_out_E_noc1_yummy;
wire tile_4_2_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_4_2_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_4_2_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_4_2_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_4_2_out_W_noc2_data;
wire tile_4_2_out_N_noc2_valid;
wire tile_4_2_out_S_noc2_valid;
wire tile_4_2_out_E_noc2_valid;
wire tile_4_2_out_W_noc2_valid;
wire tile_4_2_out_N_noc2_yummy;
wire tile_4_2_out_S_noc2_yummy;
wire tile_4_2_out_E_noc2_yummy;
wire tile_4_2_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_4_2_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_4_2_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_4_2_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_4_2_out_W_noc3_data;
wire tile_4_2_out_N_noc3_valid;
wire tile_4_2_out_S_noc3_valid;
wire tile_4_2_out_E_noc3_valid;
wire tile_4_2_out_W_noc3_valid;
wire tile_4_2_out_N_noc3_yummy;
wire tile_4_2_out_S_noc3_yummy;
wire tile_4_2_out_E_noc3_yummy;
wire tile_4_2_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_5_2_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_5_2_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_5_2_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_5_2_out_W_noc1_data;
wire tile_5_2_out_N_noc1_valid;
wire tile_5_2_out_S_noc1_valid;
wire tile_5_2_out_E_noc1_valid;
wire tile_5_2_out_W_noc1_valid;
wire tile_5_2_out_N_noc1_yummy;
wire tile_5_2_out_S_noc1_yummy;
wire tile_5_2_out_E_noc1_yummy;
wire tile_5_2_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_5_2_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_5_2_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_5_2_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_5_2_out_W_noc2_data;
wire tile_5_2_out_N_noc2_valid;
wire tile_5_2_out_S_noc2_valid;
wire tile_5_2_out_E_noc2_valid;
wire tile_5_2_out_W_noc2_valid;
wire tile_5_2_out_N_noc2_yummy;
wire tile_5_2_out_S_noc2_yummy;
wire tile_5_2_out_E_noc2_yummy;
wire tile_5_2_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_5_2_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_5_2_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_5_2_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_5_2_out_W_noc3_data;
wire tile_5_2_out_N_noc3_valid;
wire tile_5_2_out_S_noc3_valid;
wire tile_5_2_out_E_noc3_valid;
wire tile_5_2_out_W_noc3_valid;
wire tile_5_2_out_N_noc3_yummy;
wire tile_5_2_out_S_noc3_yummy;
wire tile_5_2_out_E_noc3_yummy;
wire tile_5_2_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_6_2_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_6_2_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_6_2_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_6_2_out_W_noc1_data;
wire tile_6_2_out_N_noc1_valid;
wire tile_6_2_out_S_noc1_valid;
wire tile_6_2_out_E_noc1_valid;
wire tile_6_2_out_W_noc1_valid;
wire tile_6_2_out_N_noc1_yummy;
wire tile_6_2_out_S_noc1_yummy;
wire tile_6_2_out_E_noc1_yummy;
wire tile_6_2_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_6_2_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_6_2_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_6_2_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_6_2_out_W_noc2_data;
wire tile_6_2_out_N_noc2_valid;
wire tile_6_2_out_S_noc2_valid;
wire tile_6_2_out_E_noc2_valid;
wire tile_6_2_out_W_noc2_valid;
wire tile_6_2_out_N_noc2_yummy;
wire tile_6_2_out_S_noc2_yummy;
wire tile_6_2_out_E_noc2_yummy;
wire tile_6_2_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_6_2_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_6_2_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_6_2_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_6_2_out_W_noc3_data;
wire tile_6_2_out_N_noc3_valid;
wire tile_6_2_out_S_noc3_valid;
wire tile_6_2_out_E_noc3_valid;
wire tile_6_2_out_W_noc3_valid;
wire tile_6_2_out_N_noc3_yummy;
wire tile_6_2_out_S_noc3_yummy;
wire tile_6_2_out_E_noc3_yummy;
wire tile_6_2_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_7_2_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_7_2_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_7_2_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_7_2_out_W_noc1_data;
wire tile_7_2_out_N_noc1_valid;
wire tile_7_2_out_S_noc1_valid;
wire tile_7_2_out_E_noc1_valid;
wire tile_7_2_out_W_noc1_valid;
wire tile_7_2_out_N_noc1_yummy;
wire tile_7_2_out_S_noc1_yummy;
wire tile_7_2_out_E_noc1_yummy;
wire tile_7_2_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_7_2_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_7_2_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_7_2_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_7_2_out_W_noc2_data;
wire tile_7_2_out_N_noc2_valid;
wire tile_7_2_out_S_noc2_valid;
wire tile_7_2_out_E_noc2_valid;
wire tile_7_2_out_W_noc2_valid;
wire tile_7_2_out_N_noc2_yummy;
wire tile_7_2_out_S_noc2_yummy;
wire tile_7_2_out_E_noc2_yummy;
wire tile_7_2_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_7_2_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_7_2_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_7_2_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_7_2_out_W_noc3_data;
wire tile_7_2_out_N_noc3_valid;
wire tile_7_2_out_S_noc3_valid;
wire tile_7_2_out_E_noc3_valid;
wire tile_7_2_out_W_noc3_valid;
wire tile_7_2_out_N_noc3_yummy;
wire tile_7_2_out_S_noc3_yummy;
wire tile_7_2_out_E_noc3_yummy;
wire tile_7_2_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_8_2_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_8_2_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_8_2_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_8_2_out_W_noc1_data;
wire tile_8_2_out_N_noc1_valid;
wire tile_8_2_out_S_noc1_valid;
wire tile_8_2_out_E_noc1_valid;
wire tile_8_2_out_W_noc1_valid;
wire tile_8_2_out_N_noc1_yummy;
wire tile_8_2_out_S_noc1_yummy;
wire tile_8_2_out_E_noc1_yummy;
wire tile_8_2_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_8_2_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_8_2_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_8_2_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_8_2_out_W_noc2_data;
wire tile_8_2_out_N_noc2_valid;
wire tile_8_2_out_S_noc2_valid;
wire tile_8_2_out_E_noc2_valid;
wire tile_8_2_out_W_noc2_valid;
wire tile_8_2_out_N_noc2_yummy;
wire tile_8_2_out_S_noc2_yummy;
wire tile_8_2_out_E_noc2_yummy;
wire tile_8_2_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_8_2_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_8_2_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_8_2_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_8_2_out_W_noc3_data;
wire tile_8_2_out_N_noc3_valid;
wire tile_8_2_out_S_noc3_valid;
wire tile_8_2_out_E_noc3_valid;
wire tile_8_2_out_W_noc3_valid;
wire tile_8_2_out_N_noc3_yummy;
wire tile_8_2_out_S_noc3_yummy;
wire tile_8_2_out_E_noc3_yummy;
wire tile_8_2_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_9_2_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_9_2_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_9_2_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_9_2_out_W_noc1_data;
wire tile_9_2_out_N_noc1_valid;
wire tile_9_2_out_S_noc1_valid;
wire tile_9_2_out_E_noc1_valid;
wire tile_9_2_out_W_noc1_valid;
wire tile_9_2_out_N_noc1_yummy;
wire tile_9_2_out_S_noc1_yummy;
wire tile_9_2_out_E_noc1_yummy;
wire tile_9_2_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_9_2_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_9_2_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_9_2_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_9_2_out_W_noc2_data;
wire tile_9_2_out_N_noc2_valid;
wire tile_9_2_out_S_noc2_valid;
wire tile_9_2_out_E_noc2_valid;
wire tile_9_2_out_W_noc2_valid;
wire tile_9_2_out_N_noc2_yummy;
wire tile_9_2_out_S_noc2_yummy;
wire tile_9_2_out_E_noc2_yummy;
wire tile_9_2_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_9_2_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_9_2_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_9_2_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_9_2_out_W_noc3_data;
wire tile_9_2_out_N_noc3_valid;
wire tile_9_2_out_S_noc3_valid;
wire tile_9_2_out_E_noc3_valid;
wire tile_9_2_out_W_noc3_valid;
wire tile_9_2_out_N_noc3_yummy;
wire tile_9_2_out_S_noc3_yummy;
wire tile_9_2_out_E_noc3_yummy;
wire tile_9_2_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_10_2_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_10_2_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_10_2_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_10_2_out_W_noc1_data;
wire tile_10_2_out_N_noc1_valid;
wire tile_10_2_out_S_noc1_valid;
wire tile_10_2_out_E_noc1_valid;
wire tile_10_2_out_W_noc1_valid;
wire tile_10_2_out_N_noc1_yummy;
wire tile_10_2_out_S_noc1_yummy;
wire tile_10_2_out_E_noc1_yummy;
wire tile_10_2_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_10_2_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_10_2_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_10_2_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_10_2_out_W_noc2_data;
wire tile_10_2_out_N_noc2_valid;
wire tile_10_2_out_S_noc2_valid;
wire tile_10_2_out_E_noc2_valid;
wire tile_10_2_out_W_noc2_valid;
wire tile_10_2_out_N_noc2_yummy;
wire tile_10_2_out_S_noc2_yummy;
wire tile_10_2_out_E_noc2_yummy;
wire tile_10_2_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_10_2_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_10_2_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_10_2_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_10_2_out_W_noc3_data;
wire tile_10_2_out_N_noc3_valid;
wire tile_10_2_out_S_noc3_valid;
wire tile_10_2_out_E_noc3_valid;
wire tile_10_2_out_W_noc3_valid;
wire tile_10_2_out_N_noc3_yummy;
wire tile_10_2_out_S_noc3_yummy;
wire tile_10_2_out_E_noc3_yummy;
wire tile_10_2_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_11_2_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_11_2_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_11_2_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_11_2_out_W_noc1_data;
wire tile_11_2_out_N_noc1_valid;
wire tile_11_2_out_S_noc1_valid;
wire tile_11_2_out_E_noc1_valid;
wire tile_11_2_out_W_noc1_valid;
wire tile_11_2_out_N_noc1_yummy;
wire tile_11_2_out_S_noc1_yummy;
wire tile_11_2_out_E_noc1_yummy;
wire tile_11_2_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_11_2_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_11_2_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_11_2_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_11_2_out_W_noc2_data;
wire tile_11_2_out_N_noc2_valid;
wire tile_11_2_out_S_noc2_valid;
wire tile_11_2_out_E_noc2_valid;
wire tile_11_2_out_W_noc2_valid;
wire tile_11_2_out_N_noc2_yummy;
wire tile_11_2_out_S_noc2_yummy;
wire tile_11_2_out_E_noc2_yummy;
wire tile_11_2_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_11_2_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_11_2_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_11_2_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_11_2_out_W_noc3_data;
wire tile_11_2_out_N_noc3_valid;
wire tile_11_2_out_S_noc3_valid;
wire tile_11_2_out_E_noc3_valid;
wire tile_11_2_out_W_noc3_valid;
wire tile_11_2_out_N_noc3_yummy;
wire tile_11_2_out_S_noc3_yummy;
wire tile_11_2_out_E_noc3_yummy;
wire tile_11_2_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_12_2_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_12_2_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_12_2_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_12_2_out_W_noc1_data;
wire tile_12_2_out_N_noc1_valid;
wire tile_12_2_out_S_noc1_valid;
wire tile_12_2_out_E_noc1_valid;
wire tile_12_2_out_W_noc1_valid;
wire tile_12_2_out_N_noc1_yummy;
wire tile_12_2_out_S_noc1_yummy;
wire tile_12_2_out_E_noc1_yummy;
wire tile_12_2_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_12_2_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_12_2_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_12_2_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_12_2_out_W_noc2_data;
wire tile_12_2_out_N_noc2_valid;
wire tile_12_2_out_S_noc2_valid;
wire tile_12_2_out_E_noc2_valid;
wire tile_12_2_out_W_noc2_valid;
wire tile_12_2_out_N_noc2_yummy;
wire tile_12_2_out_S_noc2_yummy;
wire tile_12_2_out_E_noc2_yummy;
wire tile_12_2_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_12_2_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_12_2_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_12_2_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_12_2_out_W_noc3_data;
wire tile_12_2_out_N_noc3_valid;
wire tile_12_2_out_S_noc3_valid;
wire tile_12_2_out_E_noc3_valid;
wire tile_12_2_out_W_noc3_valid;
wire tile_12_2_out_N_noc3_yummy;
wire tile_12_2_out_S_noc3_yummy;
wire tile_12_2_out_E_noc3_yummy;
wire tile_12_2_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_13_2_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_13_2_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_13_2_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_13_2_out_W_noc1_data;
wire tile_13_2_out_N_noc1_valid;
wire tile_13_2_out_S_noc1_valid;
wire tile_13_2_out_E_noc1_valid;
wire tile_13_2_out_W_noc1_valid;
wire tile_13_2_out_N_noc1_yummy;
wire tile_13_2_out_S_noc1_yummy;
wire tile_13_2_out_E_noc1_yummy;
wire tile_13_2_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_13_2_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_13_2_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_13_2_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_13_2_out_W_noc2_data;
wire tile_13_2_out_N_noc2_valid;
wire tile_13_2_out_S_noc2_valid;
wire tile_13_2_out_E_noc2_valid;
wire tile_13_2_out_W_noc2_valid;
wire tile_13_2_out_N_noc2_yummy;
wire tile_13_2_out_S_noc2_yummy;
wire tile_13_2_out_E_noc2_yummy;
wire tile_13_2_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_13_2_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_13_2_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_13_2_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_13_2_out_W_noc3_data;
wire tile_13_2_out_N_noc3_valid;
wire tile_13_2_out_S_noc3_valid;
wire tile_13_2_out_E_noc3_valid;
wire tile_13_2_out_W_noc3_valid;
wire tile_13_2_out_N_noc3_yummy;
wire tile_13_2_out_S_noc3_yummy;
wire tile_13_2_out_E_noc3_yummy;
wire tile_13_2_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_14_2_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_14_2_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_14_2_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_14_2_out_W_noc1_data;
wire tile_14_2_out_N_noc1_valid;
wire tile_14_2_out_S_noc1_valid;
wire tile_14_2_out_E_noc1_valid;
wire tile_14_2_out_W_noc1_valid;
wire tile_14_2_out_N_noc1_yummy;
wire tile_14_2_out_S_noc1_yummy;
wire tile_14_2_out_E_noc1_yummy;
wire tile_14_2_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_14_2_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_14_2_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_14_2_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_14_2_out_W_noc2_data;
wire tile_14_2_out_N_noc2_valid;
wire tile_14_2_out_S_noc2_valid;
wire tile_14_2_out_E_noc2_valid;
wire tile_14_2_out_W_noc2_valid;
wire tile_14_2_out_N_noc2_yummy;
wire tile_14_2_out_S_noc2_yummy;
wire tile_14_2_out_E_noc2_yummy;
wire tile_14_2_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_14_2_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_14_2_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_14_2_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_14_2_out_W_noc3_data;
wire tile_14_2_out_N_noc3_valid;
wire tile_14_2_out_S_noc3_valid;
wire tile_14_2_out_E_noc3_valid;
wire tile_14_2_out_W_noc3_valid;
wire tile_14_2_out_N_noc3_yummy;
wire tile_14_2_out_S_noc3_yummy;
wire tile_14_2_out_E_noc3_yummy;
wire tile_14_2_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_15_2_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_15_2_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_15_2_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_15_2_out_W_noc1_data;
wire tile_15_2_out_N_noc1_valid;
wire tile_15_2_out_S_noc1_valid;
wire tile_15_2_out_E_noc1_valid;
wire tile_15_2_out_W_noc1_valid;
wire tile_15_2_out_N_noc1_yummy;
wire tile_15_2_out_S_noc1_yummy;
wire tile_15_2_out_E_noc1_yummy;
wire tile_15_2_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_15_2_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_15_2_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_15_2_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_15_2_out_W_noc2_data;
wire tile_15_2_out_N_noc2_valid;
wire tile_15_2_out_S_noc2_valid;
wire tile_15_2_out_E_noc2_valid;
wire tile_15_2_out_W_noc2_valid;
wire tile_15_2_out_N_noc2_yummy;
wire tile_15_2_out_S_noc2_yummy;
wire tile_15_2_out_E_noc2_yummy;
wire tile_15_2_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_15_2_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_15_2_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_15_2_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_15_2_out_W_noc3_data;
wire tile_15_2_out_N_noc3_valid;
wire tile_15_2_out_S_noc3_valid;
wire tile_15_2_out_E_noc3_valid;
wire tile_15_2_out_W_noc3_valid;
wire tile_15_2_out_N_noc3_yummy;
wire tile_15_2_out_S_noc3_yummy;
wire tile_15_2_out_E_noc3_yummy;
wire tile_15_2_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_0_3_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_0_3_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_0_3_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_0_3_out_W_noc1_data;
wire tile_0_3_out_N_noc1_valid;
wire tile_0_3_out_S_noc1_valid;
wire tile_0_3_out_E_noc1_valid;
wire tile_0_3_out_W_noc1_valid;
wire tile_0_3_out_N_noc1_yummy;
wire tile_0_3_out_S_noc1_yummy;
wire tile_0_3_out_E_noc1_yummy;
wire tile_0_3_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_0_3_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_0_3_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_0_3_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_0_3_out_W_noc2_data;
wire tile_0_3_out_N_noc2_valid;
wire tile_0_3_out_S_noc2_valid;
wire tile_0_3_out_E_noc2_valid;
wire tile_0_3_out_W_noc2_valid;
wire tile_0_3_out_N_noc2_yummy;
wire tile_0_3_out_S_noc2_yummy;
wire tile_0_3_out_E_noc2_yummy;
wire tile_0_3_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_0_3_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_0_3_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_0_3_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_0_3_out_W_noc3_data;
wire tile_0_3_out_N_noc3_valid;
wire tile_0_3_out_S_noc3_valid;
wire tile_0_3_out_E_noc3_valid;
wire tile_0_3_out_W_noc3_valid;
wire tile_0_3_out_N_noc3_yummy;
wire tile_0_3_out_S_noc3_yummy;
wire tile_0_3_out_E_noc3_yummy;
wire tile_0_3_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_1_3_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_1_3_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_1_3_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_1_3_out_W_noc1_data;
wire tile_1_3_out_N_noc1_valid;
wire tile_1_3_out_S_noc1_valid;
wire tile_1_3_out_E_noc1_valid;
wire tile_1_3_out_W_noc1_valid;
wire tile_1_3_out_N_noc1_yummy;
wire tile_1_3_out_S_noc1_yummy;
wire tile_1_3_out_E_noc1_yummy;
wire tile_1_3_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_1_3_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_1_3_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_1_3_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_1_3_out_W_noc2_data;
wire tile_1_3_out_N_noc2_valid;
wire tile_1_3_out_S_noc2_valid;
wire tile_1_3_out_E_noc2_valid;
wire tile_1_3_out_W_noc2_valid;
wire tile_1_3_out_N_noc2_yummy;
wire tile_1_3_out_S_noc2_yummy;
wire tile_1_3_out_E_noc2_yummy;
wire tile_1_3_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_1_3_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_1_3_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_1_3_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_1_3_out_W_noc3_data;
wire tile_1_3_out_N_noc3_valid;
wire tile_1_3_out_S_noc3_valid;
wire tile_1_3_out_E_noc3_valid;
wire tile_1_3_out_W_noc3_valid;
wire tile_1_3_out_N_noc3_yummy;
wire tile_1_3_out_S_noc3_yummy;
wire tile_1_3_out_E_noc3_yummy;
wire tile_1_3_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_2_3_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_2_3_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_2_3_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_2_3_out_W_noc1_data;
wire tile_2_3_out_N_noc1_valid;
wire tile_2_3_out_S_noc1_valid;
wire tile_2_3_out_E_noc1_valid;
wire tile_2_3_out_W_noc1_valid;
wire tile_2_3_out_N_noc1_yummy;
wire tile_2_3_out_S_noc1_yummy;
wire tile_2_3_out_E_noc1_yummy;
wire tile_2_3_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_2_3_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_2_3_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_2_3_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_2_3_out_W_noc2_data;
wire tile_2_3_out_N_noc2_valid;
wire tile_2_3_out_S_noc2_valid;
wire tile_2_3_out_E_noc2_valid;
wire tile_2_3_out_W_noc2_valid;
wire tile_2_3_out_N_noc2_yummy;
wire tile_2_3_out_S_noc2_yummy;
wire tile_2_3_out_E_noc2_yummy;
wire tile_2_3_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_2_3_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_2_3_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_2_3_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_2_3_out_W_noc3_data;
wire tile_2_3_out_N_noc3_valid;
wire tile_2_3_out_S_noc3_valid;
wire tile_2_3_out_E_noc3_valid;
wire tile_2_3_out_W_noc3_valid;
wire tile_2_3_out_N_noc3_yummy;
wire tile_2_3_out_S_noc3_yummy;
wire tile_2_3_out_E_noc3_yummy;
wire tile_2_3_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_3_3_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_3_3_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_3_3_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_3_3_out_W_noc1_data;
wire tile_3_3_out_N_noc1_valid;
wire tile_3_3_out_S_noc1_valid;
wire tile_3_3_out_E_noc1_valid;
wire tile_3_3_out_W_noc1_valid;
wire tile_3_3_out_N_noc1_yummy;
wire tile_3_3_out_S_noc1_yummy;
wire tile_3_3_out_E_noc1_yummy;
wire tile_3_3_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_3_3_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_3_3_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_3_3_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_3_3_out_W_noc2_data;
wire tile_3_3_out_N_noc2_valid;
wire tile_3_3_out_S_noc2_valid;
wire tile_3_3_out_E_noc2_valid;
wire tile_3_3_out_W_noc2_valid;
wire tile_3_3_out_N_noc2_yummy;
wire tile_3_3_out_S_noc2_yummy;
wire tile_3_3_out_E_noc2_yummy;
wire tile_3_3_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_3_3_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_3_3_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_3_3_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_3_3_out_W_noc3_data;
wire tile_3_3_out_N_noc3_valid;
wire tile_3_3_out_S_noc3_valid;
wire tile_3_3_out_E_noc3_valid;
wire tile_3_3_out_W_noc3_valid;
wire tile_3_3_out_N_noc3_yummy;
wire tile_3_3_out_S_noc3_yummy;
wire tile_3_3_out_E_noc3_yummy;
wire tile_3_3_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_4_3_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_4_3_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_4_3_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_4_3_out_W_noc1_data;
wire tile_4_3_out_N_noc1_valid;
wire tile_4_3_out_S_noc1_valid;
wire tile_4_3_out_E_noc1_valid;
wire tile_4_3_out_W_noc1_valid;
wire tile_4_3_out_N_noc1_yummy;
wire tile_4_3_out_S_noc1_yummy;
wire tile_4_3_out_E_noc1_yummy;
wire tile_4_3_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_4_3_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_4_3_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_4_3_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_4_3_out_W_noc2_data;
wire tile_4_3_out_N_noc2_valid;
wire tile_4_3_out_S_noc2_valid;
wire tile_4_3_out_E_noc2_valid;
wire tile_4_3_out_W_noc2_valid;
wire tile_4_3_out_N_noc2_yummy;
wire tile_4_3_out_S_noc2_yummy;
wire tile_4_3_out_E_noc2_yummy;
wire tile_4_3_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_4_3_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_4_3_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_4_3_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_4_3_out_W_noc3_data;
wire tile_4_3_out_N_noc3_valid;
wire tile_4_3_out_S_noc3_valid;
wire tile_4_3_out_E_noc3_valid;
wire tile_4_3_out_W_noc3_valid;
wire tile_4_3_out_N_noc3_yummy;
wire tile_4_3_out_S_noc3_yummy;
wire tile_4_3_out_E_noc3_yummy;
wire tile_4_3_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_5_3_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_5_3_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_5_3_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_5_3_out_W_noc1_data;
wire tile_5_3_out_N_noc1_valid;
wire tile_5_3_out_S_noc1_valid;
wire tile_5_3_out_E_noc1_valid;
wire tile_5_3_out_W_noc1_valid;
wire tile_5_3_out_N_noc1_yummy;
wire tile_5_3_out_S_noc1_yummy;
wire tile_5_3_out_E_noc1_yummy;
wire tile_5_3_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_5_3_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_5_3_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_5_3_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_5_3_out_W_noc2_data;
wire tile_5_3_out_N_noc2_valid;
wire tile_5_3_out_S_noc2_valid;
wire tile_5_3_out_E_noc2_valid;
wire tile_5_3_out_W_noc2_valid;
wire tile_5_3_out_N_noc2_yummy;
wire tile_5_3_out_S_noc2_yummy;
wire tile_5_3_out_E_noc2_yummy;
wire tile_5_3_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_5_3_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_5_3_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_5_3_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_5_3_out_W_noc3_data;
wire tile_5_3_out_N_noc3_valid;
wire tile_5_3_out_S_noc3_valid;
wire tile_5_3_out_E_noc3_valid;
wire tile_5_3_out_W_noc3_valid;
wire tile_5_3_out_N_noc3_yummy;
wire tile_5_3_out_S_noc3_yummy;
wire tile_5_3_out_E_noc3_yummy;
wire tile_5_3_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_6_3_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_6_3_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_6_3_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_6_3_out_W_noc1_data;
wire tile_6_3_out_N_noc1_valid;
wire tile_6_3_out_S_noc1_valid;
wire tile_6_3_out_E_noc1_valid;
wire tile_6_3_out_W_noc1_valid;
wire tile_6_3_out_N_noc1_yummy;
wire tile_6_3_out_S_noc1_yummy;
wire tile_6_3_out_E_noc1_yummy;
wire tile_6_3_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_6_3_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_6_3_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_6_3_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_6_3_out_W_noc2_data;
wire tile_6_3_out_N_noc2_valid;
wire tile_6_3_out_S_noc2_valid;
wire tile_6_3_out_E_noc2_valid;
wire tile_6_3_out_W_noc2_valid;
wire tile_6_3_out_N_noc2_yummy;
wire tile_6_3_out_S_noc2_yummy;
wire tile_6_3_out_E_noc2_yummy;
wire tile_6_3_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_6_3_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_6_3_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_6_3_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_6_3_out_W_noc3_data;
wire tile_6_3_out_N_noc3_valid;
wire tile_6_3_out_S_noc3_valid;
wire tile_6_3_out_E_noc3_valid;
wire tile_6_3_out_W_noc3_valid;
wire tile_6_3_out_N_noc3_yummy;
wire tile_6_3_out_S_noc3_yummy;
wire tile_6_3_out_E_noc3_yummy;
wire tile_6_3_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_7_3_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_7_3_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_7_3_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_7_3_out_W_noc1_data;
wire tile_7_3_out_N_noc1_valid;
wire tile_7_3_out_S_noc1_valid;
wire tile_7_3_out_E_noc1_valid;
wire tile_7_3_out_W_noc1_valid;
wire tile_7_3_out_N_noc1_yummy;
wire tile_7_3_out_S_noc1_yummy;
wire tile_7_3_out_E_noc1_yummy;
wire tile_7_3_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_7_3_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_7_3_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_7_3_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_7_3_out_W_noc2_data;
wire tile_7_3_out_N_noc2_valid;
wire tile_7_3_out_S_noc2_valid;
wire tile_7_3_out_E_noc2_valid;
wire tile_7_3_out_W_noc2_valid;
wire tile_7_3_out_N_noc2_yummy;
wire tile_7_3_out_S_noc2_yummy;
wire tile_7_3_out_E_noc2_yummy;
wire tile_7_3_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_7_3_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_7_3_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_7_3_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_7_3_out_W_noc3_data;
wire tile_7_3_out_N_noc3_valid;
wire tile_7_3_out_S_noc3_valid;
wire tile_7_3_out_E_noc3_valid;
wire tile_7_3_out_W_noc3_valid;
wire tile_7_3_out_N_noc3_yummy;
wire tile_7_3_out_S_noc3_yummy;
wire tile_7_3_out_E_noc3_yummy;
wire tile_7_3_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_8_3_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_8_3_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_8_3_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_8_3_out_W_noc1_data;
wire tile_8_3_out_N_noc1_valid;
wire tile_8_3_out_S_noc1_valid;
wire tile_8_3_out_E_noc1_valid;
wire tile_8_3_out_W_noc1_valid;
wire tile_8_3_out_N_noc1_yummy;
wire tile_8_3_out_S_noc1_yummy;
wire tile_8_3_out_E_noc1_yummy;
wire tile_8_3_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_8_3_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_8_3_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_8_3_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_8_3_out_W_noc2_data;
wire tile_8_3_out_N_noc2_valid;
wire tile_8_3_out_S_noc2_valid;
wire tile_8_3_out_E_noc2_valid;
wire tile_8_3_out_W_noc2_valid;
wire tile_8_3_out_N_noc2_yummy;
wire tile_8_3_out_S_noc2_yummy;
wire tile_8_3_out_E_noc2_yummy;
wire tile_8_3_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_8_3_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_8_3_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_8_3_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_8_3_out_W_noc3_data;
wire tile_8_3_out_N_noc3_valid;
wire tile_8_3_out_S_noc3_valid;
wire tile_8_3_out_E_noc3_valid;
wire tile_8_3_out_W_noc3_valid;
wire tile_8_3_out_N_noc3_yummy;
wire tile_8_3_out_S_noc3_yummy;
wire tile_8_3_out_E_noc3_yummy;
wire tile_8_3_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_9_3_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_9_3_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_9_3_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_9_3_out_W_noc1_data;
wire tile_9_3_out_N_noc1_valid;
wire tile_9_3_out_S_noc1_valid;
wire tile_9_3_out_E_noc1_valid;
wire tile_9_3_out_W_noc1_valid;
wire tile_9_3_out_N_noc1_yummy;
wire tile_9_3_out_S_noc1_yummy;
wire tile_9_3_out_E_noc1_yummy;
wire tile_9_3_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_9_3_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_9_3_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_9_3_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_9_3_out_W_noc2_data;
wire tile_9_3_out_N_noc2_valid;
wire tile_9_3_out_S_noc2_valid;
wire tile_9_3_out_E_noc2_valid;
wire tile_9_3_out_W_noc2_valid;
wire tile_9_3_out_N_noc2_yummy;
wire tile_9_3_out_S_noc2_yummy;
wire tile_9_3_out_E_noc2_yummy;
wire tile_9_3_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_9_3_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_9_3_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_9_3_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_9_3_out_W_noc3_data;
wire tile_9_3_out_N_noc3_valid;
wire tile_9_3_out_S_noc3_valid;
wire tile_9_3_out_E_noc3_valid;
wire tile_9_3_out_W_noc3_valid;
wire tile_9_3_out_N_noc3_yummy;
wire tile_9_3_out_S_noc3_yummy;
wire tile_9_3_out_E_noc3_yummy;
wire tile_9_3_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_10_3_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_10_3_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_10_3_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_10_3_out_W_noc1_data;
wire tile_10_3_out_N_noc1_valid;
wire tile_10_3_out_S_noc1_valid;
wire tile_10_3_out_E_noc1_valid;
wire tile_10_3_out_W_noc1_valid;
wire tile_10_3_out_N_noc1_yummy;
wire tile_10_3_out_S_noc1_yummy;
wire tile_10_3_out_E_noc1_yummy;
wire tile_10_3_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_10_3_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_10_3_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_10_3_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_10_3_out_W_noc2_data;
wire tile_10_3_out_N_noc2_valid;
wire tile_10_3_out_S_noc2_valid;
wire tile_10_3_out_E_noc2_valid;
wire tile_10_3_out_W_noc2_valid;
wire tile_10_3_out_N_noc2_yummy;
wire tile_10_3_out_S_noc2_yummy;
wire tile_10_3_out_E_noc2_yummy;
wire tile_10_3_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_10_3_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_10_3_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_10_3_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_10_3_out_W_noc3_data;
wire tile_10_3_out_N_noc3_valid;
wire tile_10_3_out_S_noc3_valid;
wire tile_10_3_out_E_noc3_valid;
wire tile_10_3_out_W_noc3_valid;
wire tile_10_3_out_N_noc3_yummy;
wire tile_10_3_out_S_noc3_yummy;
wire tile_10_3_out_E_noc3_yummy;
wire tile_10_3_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_11_3_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_11_3_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_11_3_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_11_3_out_W_noc1_data;
wire tile_11_3_out_N_noc1_valid;
wire tile_11_3_out_S_noc1_valid;
wire tile_11_3_out_E_noc1_valid;
wire tile_11_3_out_W_noc1_valid;
wire tile_11_3_out_N_noc1_yummy;
wire tile_11_3_out_S_noc1_yummy;
wire tile_11_3_out_E_noc1_yummy;
wire tile_11_3_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_11_3_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_11_3_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_11_3_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_11_3_out_W_noc2_data;
wire tile_11_3_out_N_noc2_valid;
wire tile_11_3_out_S_noc2_valid;
wire tile_11_3_out_E_noc2_valid;
wire tile_11_3_out_W_noc2_valid;
wire tile_11_3_out_N_noc2_yummy;
wire tile_11_3_out_S_noc2_yummy;
wire tile_11_3_out_E_noc2_yummy;
wire tile_11_3_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_11_3_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_11_3_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_11_3_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_11_3_out_W_noc3_data;
wire tile_11_3_out_N_noc3_valid;
wire tile_11_3_out_S_noc3_valid;
wire tile_11_3_out_E_noc3_valid;
wire tile_11_3_out_W_noc3_valid;
wire tile_11_3_out_N_noc3_yummy;
wire tile_11_3_out_S_noc3_yummy;
wire tile_11_3_out_E_noc3_yummy;
wire tile_11_3_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_12_3_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_12_3_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_12_3_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_12_3_out_W_noc1_data;
wire tile_12_3_out_N_noc1_valid;
wire tile_12_3_out_S_noc1_valid;
wire tile_12_3_out_E_noc1_valid;
wire tile_12_3_out_W_noc1_valid;
wire tile_12_3_out_N_noc1_yummy;
wire tile_12_3_out_S_noc1_yummy;
wire tile_12_3_out_E_noc1_yummy;
wire tile_12_3_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_12_3_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_12_3_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_12_3_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_12_3_out_W_noc2_data;
wire tile_12_3_out_N_noc2_valid;
wire tile_12_3_out_S_noc2_valid;
wire tile_12_3_out_E_noc2_valid;
wire tile_12_3_out_W_noc2_valid;
wire tile_12_3_out_N_noc2_yummy;
wire tile_12_3_out_S_noc2_yummy;
wire tile_12_3_out_E_noc2_yummy;
wire tile_12_3_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_12_3_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_12_3_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_12_3_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_12_3_out_W_noc3_data;
wire tile_12_3_out_N_noc3_valid;
wire tile_12_3_out_S_noc3_valid;
wire tile_12_3_out_E_noc3_valid;
wire tile_12_3_out_W_noc3_valid;
wire tile_12_3_out_N_noc3_yummy;
wire tile_12_3_out_S_noc3_yummy;
wire tile_12_3_out_E_noc3_yummy;
wire tile_12_3_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_13_3_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_13_3_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_13_3_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_13_3_out_W_noc1_data;
wire tile_13_3_out_N_noc1_valid;
wire tile_13_3_out_S_noc1_valid;
wire tile_13_3_out_E_noc1_valid;
wire tile_13_3_out_W_noc1_valid;
wire tile_13_3_out_N_noc1_yummy;
wire tile_13_3_out_S_noc1_yummy;
wire tile_13_3_out_E_noc1_yummy;
wire tile_13_3_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_13_3_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_13_3_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_13_3_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_13_3_out_W_noc2_data;
wire tile_13_3_out_N_noc2_valid;
wire tile_13_3_out_S_noc2_valid;
wire tile_13_3_out_E_noc2_valid;
wire tile_13_3_out_W_noc2_valid;
wire tile_13_3_out_N_noc2_yummy;
wire tile_13_3_out_S_noc2_yummy;
wire tile_13_3_out_E_noc2_yummy;
wire tile_13_3_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_13_3_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_13_3_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_13_3_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_13_3_out_W_noc3_data;
wire tile_13_3_out_N_noc3_valid;
wire tile_13_3_out_S_noc3_valid;
wire tile_13_3_out_E_noc3_valid;
wire tile_13_3_out_W_noc3_valid;
wire tile_13_3_out_N_noc3_yummy;
wire tile_13_3_out_S_noc3_yummy;
wire tile_13_3_out_E_noc3_yummy;
wire tile_13_3_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_14_3_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_14_3_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_14_3_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_14_3_out_W_noc1_data;
wire tile_14_3_out_N_noc1_valid;
wire tile_14_3_out_S_noc1_valid;
wire tile_14_3_out_E_noc1_valid;
wire tile_14_3_out_W_noc1_valid;
wire tile_14_3_out_N_noc1_yummy;
wire tile_14_3_out_S_noc1_yummy;
wire tile_14_3_out_E_noc1_yummy;
wire tile_14_3_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_14_3_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_14_3_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_14_3_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_14_3_out_W_noc2_data;
wire tile_14_3_out_N_noc2_valid;
wire tile_14_3_out_S_noc2_valid;
wire tile_14_3_out_E_noc2_valid;
wire tile_14_3_out_W_noc2_valid;
wire tile_14_3_out_N_noc2_yummy;
wire tile_14_3_out_S_noc2_yummy;
wire tile_14_3_out_E_noc2_yummy;
wire tile_14_3_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_14_3_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_14_3_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_14_3_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_14_3_out_W_noc3_data;
wire tile_14_3_out_N_noc3_valid;
wire tile_14_3_out_S_noc3_valid;
wire tile_14_3_out_E_noc3_valid;
wire tile_14_3_out_W_noc3_valid;
wire tile_14_3_out_N_noc3_yummy;
wire tile_14_3_out_S_noc3_yummy;
wire tile_14_3_out_E_noc3_yummy;
wire tile_14_3_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_15_3_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_15_3_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_15_3_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_15_3_out_W_noc1_data;
wire tile_15_3_out_N_noc1_valid;
wire tile_15_3_out_S_noc1_valid;
wire tile_15_3_out_E_noc1_valid;
wire tile_15_3_out_W_noc1_valid;
wire tile_15_3_out_N_noc1_yummy;
wire tile_15_3_out_S_noc1_yummy;
wire tile_15_3_out_E_noc1_yummy;
wire tile_15_3_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_15_3_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_15_3_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_15_3_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_15_3_out_W_noc2_data;
wire tile_15_3_out_N_noc2_valid;
wire tile_15_3_out_S_noc2_valid;
wire tile_15_3_out_E_noc2_valid;
wire tile_15_3_out_W_noc2_valid;
wire tile_15_3_out_N_noc2_yummy;
wire tile_15_3_out_S_noc2_yummy;
wire tile_15_3_out_E_noc2_yummy;
wire tile_15_3_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_15_3_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_15_3_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_15_3_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_15_3_out_W_noc3_data;
wire tile_15_3_out_N_noc3_valid;
wire tile_15_3_out_S_noc3_valid;
wire tile_15_3_out_E_noc3_valid;
wire tile_15_3_out_W_noc3_valid;
wire tile_15_3_out_N_noc3_yummy;
wire tile_15_3_out_S_noc3_yummy;
wire tile_15_3_out_E_noc3_yummy;
wire tile_15_3_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_0_4_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_0_4_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_0_4_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_0_4_out_W_noc1_data;
wire tile_0_4_out_N_noc1_valid;
wire tile_0_4_out_S_noc1_valid;
wire tile_0_4_out_E_noc1_valid;
wire tile_0_4_out_W_noc1_valid;
wire tile_0_4_out_N_noc1_yummy;
wire tile_0_4_out_S_noc1_yummy;
wire tile_0_4_out_E_noc1_yummy;
wire tile_0_4_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_0_4_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_0_4_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_0_4_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_0_4_out_W_noc2_data;
wire tile_0_4_out_N_noc2_valid;
wire tile_0_4_out_S_noc2_valid;
wire tile_0_4_out_E_noc2_valid;
wire tile_0_4_out_W_noc2_valid;
wire tile_0_4_out_N_noc2_yummy;
wire tile_0_4_out_S_noc2_yummy;
wire tile_0_4_out_E_noc2_yummy;
wire tile_0_4_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_0_4_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_0_4_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_0_4_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_0_4_out_W_noc3_data;
wire tile_0_4_out_N_noc3_valid;
wire tile_0_4_out_S_noc3_valid;
wire tile_0_4_out_E_noc3_valid;
wire tile_0_4_out_W_noc3_valid;
wire tile_0_4_out_N_noc3_yummy;
wire tile_0_4_out_S_noc3_yummy;
wire tile_0_4_out_E_noc3_yummy;
wire tile_0_4_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_1_4_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_1_4_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_1_4_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_1_4_out_W_noc1_data;
wire tile_1_4_out_N_noc1_valid;
wire tile_1_4_out_S_noc1_valid;
wire tile_1_4_out_E_noc1_valid;
wire tile_1_4_out_W_noc1_valid;
wire tile_1_4_out_N_noc1_yummy;
wire tile_1_4_out_S_noc1_yummy;
wire tile_1_4_out_E_noc1_yummy;
wire tile_1_4_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_1_4_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_1_4_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_1_4_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_1_4_out_W_noc2_data;
wire tile_1_4_out_N_noc2_valid;
wire tile_1_4_out_S_noc2_valid;
wire tile_1_4_out_E_noc2_valid;
wire tile_1_4_out_W_noc2_valid;
wire tile_1_4_out_N_noc2_yummy;
wire tile_1_4_out_S_noc2_yummy;
wire tile_1_4_out_E_noc2_yummy;
wire tile_1_4_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_1_4_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_1_4_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_1_4_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_1_4_out_W_noc3_data;
wire tile_1_4_out_N_noc3_valid;
wire tile_1_4_out_S_noc3_valid;
wire tile_1_4_out_E_noc3_valid;
wire tile_1_4_out_W_noc3_valid;
wire tile_1_4_out_N_noc3_yummy;
wire tile_1_4_out_S_noc3_yummy;
wire tile_1_4_out_E_noc3_yummy;
wire tile_1_4_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_2_4_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_2_4_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_2_4_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_2_4_out_W_noc1_data;
wire tile_2_4_out_N_noc1_valid;
wire tile_2_4_out_S_noc1_valid;
wire tile_2_4_out_E_noc1_valid;
wire tile_2_4_out_W_noc1_valid;
wire tile_2_4_out_N_noc1_yummy;
wire tile_2_4_out_S_noc1_yummy;
wire tile_2_4_out_E_noc1_yummy;
wire tile_2_4_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_2_4_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_2_4_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_2_4_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_2_4_out_W_noc2_data;
wire tile_2_4_out_N_noc2_valid;
wire tile_2_4_out_S_noc2_valid;
wire tile_2_4_out_E_noc2_valid;
wire tile_2_4_out_W_noc2_valid;
wire tile_2_4_out_N_noc2_yummy;
wire tile_2_4_out_S_noc2_yummy;
wire tile_2_4_out_E_noc2_yummy;
wire tile_2_4_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_2_4_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_2_4_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_2_4_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_2_4_out_W_noc3_data;
wire tile_2_4_out_N_noc3_valid;
wire tile_2_4_out_S_noc3_valid;
wire tile_2_4_out_E_noc3_valid;
wire tile_2_4_out_W_noc3_valid;
wire tile_2_4_out_N_noc3_yummy;
wire tile_2_4_out_S_noc3_yummy;
wire tile_2_4_out_E_noc3_yummy;
wire tile_2_4_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_3_4_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_3_4_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_3_4_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_3_4_out_W_noc1_data;
wire tile_3_4_out_N_noc1_valid;
wire tile_3_4_out_S_noc1_valid;
wire tile_3_4_out_E_noc1_valid;
wire tile_3_4_out_W_noc1_valid;
wire tile_3_4_out_N_noc1_yummy;
wire tile_3_4_out_S_noc1_yummy;
wire tile_3_4_out_E_noc1_yummy;
wire tile_3_4_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_3_4_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_3_4_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_3_4_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_3_4_out_W_noc2_data;
wire tile_3_4_out_N_noc2_valid;
wire tile_3_4_out_S_noc2_valid;
wire tile_3_4_out_E_noc2_valid;
wire tile_3_4_out_W_noc2_valid;
wire tile_3_4_out_N_noc2_yummy;
wire tile_3_4_out_S_noc2_yummy;
wire tile_3_4_out_E_noc2_yummy;
wire tile_3_4_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_3_4_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_3_4_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_3_4_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_3_4_out_W_noc3_data;
wire tile_3_4_out_N_noc3_valid;
wire tile_3_4_out_S_noc3_valid;
wire tile_3_4_out_E_noc3_valid;
wire tile_3_4_out_W_noc3_valid;
wire tile_3_4_out_N_noc3_yummy;
wire tile_3_4_out_S_noc3_yummy;
wire tile_3_4_out_E_noc3_yummy;
wire tile_3_4_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_4_4_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_4_4_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_4_4_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_4_4_out_W_noc1_data;
wire tile_4_4_out_N_noc1_valid;
wire tile_4_4_out_S_noc1_valid;
wire tile_4_4_out_E_noc1_valid;
wire tile_4_4_out_W_noc1_valid;
wire tile_4_4_out_N_noc1_yummy;
wire tile_4_4_out_S_noc1_yummy;
wire tile_4_4_out_E_noc1_yummy;
wire tile_4_4_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_4_4_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_4_4_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_4_4_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_4_4_out_W_noc2_data;
wire tile_4_4_out_N_noc2_valid;
wire tile_4_4_out_S_noc2_valid;
wire tile_4_4_out_E_noc2_valid;
wire tile_4_4_out_W_noc2_valid;
wire tile_4_4_out_N_noc2_yummy;
wire tile_4_4_out_S_noc2_yummy;
wire tile_4_4_out_E_noc2_yummy;
wire tile_4_4_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_4_4_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_4_4_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_4_4_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_4_4_out_W_noc3_data;
wire tile_4_4_out_N_noc3_valid;
wire tile_4_4_out_S_noc3_valid;
wire tile_4_4_out_E_noc3_valid;
wire tile_4_4_out_W_noc3_valid;
wire tile_4_4_out_N_noc3_yummy;
wire tile_4_4_out_S_noc3_yummy;
wire tile_4_4_out_E_noc3_yummy;
wire tile_4_4_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_5_4_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_5_4_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_5_4_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_5_4_out_W_noc1_data;
wire tile_5_4_out_N_noc1_valid;
wire tile_5_4_out_S_noc1_valid;
wire tile_5_4_out_E_noc1_valid;
wire tile_5_4_out_W_noc1_valid;
wire tile_5_4_out_N_noc1_yummy;
wire tile_5_4_out_S_noc1_yummy;
wire tile_5_4_out_E_noc1_yummy;
wire tile_5_4_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_5_4_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_5_4_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_5_4_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_5_4_out_W_noc2_data;
wire tile_5_4_out_N_noc2_valid;
wire tile_5_4_out_S_noc2_valid;
wire tile_5_4_out_E_noc2_valid;
wire tile_5_4_out_W_noc2_valid;
wire tile_5_4_out_N_noc2_yummy;
wire tile_5_4_out_S_noc2_yummy;
wire tile_5_4_out_E_noc2_yummy;
wire tile_5_4_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_5_4_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_5_4_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_5_4_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_5_4_out_W_noc3_data;
wire tile_5_4_out_N_noc3_valid;
wire tile_5_4_out_S_noc3_valid;
wire tile_5_4_out_E_noc3_valid;
wire tile_5_4_out_W_noc3_valid;
wire tile_5_4_out_N_noc3_yummy;
wire tile_5_4_out_S_noc3_yummy;
wire tile_5_4_out_E_noc3_yummy;
wire tile_5_4_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_6_4_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_6_4_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_6_4_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_6_4_out_W_noc1_data;
wire tile_6_4_out_N_noc1_valid;
wire tile_6_4_out_S_noc1_valid;
wire tile_6_4_out_E_noc1_valid;
wire tile_6_4_out_W_noc1_valid;
wire tile_6_4_out_N_noc1_yummy;
wire tile_6_4_out_S_noc1_yummy;
wire tile_6_4_out_E_noc1_yummy;
wire tile_6_4_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_6_4_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_6_4_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_6_4_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_6_4_out_W_noc2_data;
wire tile_6_4_out_N_noc2_valid;
wire tile_6_4_out_S_noc2_valid;
wire tile_6_4_out_E_noc2_valid;
wire tile_6_4_out_W_noc2_valid;
wire tile_6_4_out_N_noc2_yummy;
wire tile_6_4_out_S_noc2_yummy;
wire tile_6_4_out_E_noc2_yummy;
wire tile_6_4_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_6_4_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_6_4_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_6_4_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_6_4_out_W_noc3_data;
wire tile_6_4_out_N_noc3_valid;
wire tile_6_4_out_S_noc3_valid;
wire tile_6_4_out_E_noc3_valid;
wire tile_6_4_out_W_noc3_valid;
wire tile_6_4_out_N_noc3_yummy;
wire tile_6_4_out_S_noc3_yummy;
wire tile_6_4_out_E_noc3_yummy;
wire tile_6_4_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_7_4_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_7_4_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_7_4_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_7_4_out_W_noc1_data;
wire tile_7_4_out_N_noc1_valid;
wire tile_7_4_out_S_noc1_valid;
wire tile_7_4_out_E_noc1_valid;
wire tile_7_4_out_W_noc1_valid;
wire tile_7_4_out_N_noc1_yummy;
wire tile_7_4_out_S_noc1_yummy;
wire tile_7_4_out_E_noc1_yummy;
wire tile_7_4_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_7_4_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_7_4_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_7_4_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_7_4_out_W_noc2_data;
wire tile_7_4_out_N_noc2_valid;
wire tile_7_4_out_S_noc2_valid;
wire tile_7_4_out_E_noc2_valid;
wire tile_7_4_out_W_noc2_valid;
wire tile_7_4_out_N_noc2_yummy;
wire tile_7_4_out_S_noc2_yummy;
wire tile_7_4_out_E_noc2_yummy;
wire tile_7_4_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_7_4_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_7_4_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_7_4_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_7_4_out_W_noc3_data;
wire tile_7_4_out_N_noc3_valid;
wire tile_7_4_out_S_noc3_valid;
wire tile_7_4_out_E_noc3_valid;
wire tile_7_4_out_W_noc3_valid;
wire tile_7_4_out_N_noc3_yummy;
wire tile_7_4_out_S_noc3_yummy;
wire tile_7_4_out_E_noc3_yummy;
wire tile_7_4_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_8_4_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_8_4_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_8_4_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_8_4_out_W_noc1_data;
wire tile_8_4_out_N_noc1_valid;
wire tile_8_4_out_S_noc1_valid;
wire tile_8_4_out_E_noc1_valid;
wire tile_8_4_out_W_noc1_valid;
wire tile_8_4_out_N_noc1_yummy;
wire tile_8_4_out_S_noc1_yummy;
wire tile_8_4_out_E_noc1_yummy;
wire tile_8_4_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_8_4_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_8_4_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_8_4_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_8_4_out_W_noc2_data;
wire tile_8_4_out_N_noc2_valid;
wire tile_8_4_out_S_noc2_valid;
wire tile_8_4_out_E_noc2_valid;
wire tile_8_4_out_W_noc2_valid;
wire tile_8_4_out_N_noc2_yummy;
wire tile_8_4_out_S_noc2_yummy;
wire tile_8_4_out_E_noc2_yummy;
wire tile_8_4_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_8_4_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_8_4_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_8_4_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_8_4_out_W_noc3_data;
wire tile_8_4_out_N_noc3_valid;
wire tile_8_4_out_S_noc3_valid;
wire tile_8_4_out_E_noc3_valid;
wire tile_8_4_out_W_noc3_valid;
wire tile_8_4_out_N_noc3_yummy;
wire tile_8_4_out_S_noc3_yummy;
wire tile_8_4_out_E_noc3_yummy;
wire tile_8_4_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_9_4_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_9_4_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_9_4_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_9_4_out_W_noc1_data;
wire tile_9_4_out_N_noc1_valid;
wire tile_9_4_out_S_noc1_valid;
wire tile_9_4_out_E_noc1_valid;
wire tile_9_4_out_W_noc1_valid;
wire tile_9_4_out_N_noc1_yummy;
wire tile_9_4_out_S_noc1_yummy;
wire tile_9_4_out_E_noc1_yummy;
wire tile_9_4_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_9_4_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_9_4_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_9_4_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_9_4_out_W_noc2_data;
wire tile_9_4_out_N_noc2_valid;
wire tile_9_4_out_S_noc2_valid;
wire tile_9_4_out_E_noc2_valid;
wire tile_9_4_out_W_noc2_valid;
wire tile_9_4_out_N_noc2_yummy;
wire tile_9_4_out_S_noc2_yummy;
wire tile_9_4_out_E_noc2_yummy;
wire tile_9_4_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_9_4_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_9_4_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_9_4_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_9_4_out_W_noc3_data;
wire tile_9_4_out_N_noc3_valid;
wire tile_9_4_out_S_noc3_valid;
wire tile_9_4_out_E_noc3_valid;
wire tile_9_4_out_W_noc3_valid;
wire tile_9_4_out_N_noc3_yummy;
wire tile_9_4_out_S_noc3_yummy;
wire tile_9_4_out_E_noc3_yummy;
wire tile_9_4_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_10_4_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_10_4_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_10_4_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_10_4_out_W_noc1_data;
wire tile_10_4_out_N_noc1_valid;
wire tile_10_4_out_S_noc1_valid;
wire tile_10_4_out_E_noc1_valid;
wire tile_10_4_out_W_noc1_valid;
wire tile_10_4_out_N_noc1_yummy;
wire tile_10_4_out_S_noc1_yummy;
wire tile_10_4_out_E_noc1_yummy;
wire tile_10_4_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_10_4_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_10_4_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_10_4_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_10_4_out_W_noc2_data;
wire tile_10_4_out_N_noc2_valid;
wire tile_10_4_out_S_noc2_valid;
wire tile_10_4_out_E_noc2_valid;
wire tile_10_4_out_W_noc2_valid;
wire tile_10_4_out_N_noc2_yummy;
wire tile_10_4_out_S_noc2_yummy;
wire tile_10_4_out_E_noc2_yummy;
wire tile_10_4_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_10_4_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_10_4_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_10_4_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_10_4_out_W_noc3_data;
wire tile_10_4_out_N_noc3_valid;
wire tile_10_4_out_S_noc3_valid;
wire tile_10_4_out_E_noc3_valid;
wire tile_10_4_out_W_noc3_valid;
wire tile_10_4_out_N_noc3_yummy;
wire tile_10_4_out_S_noc3_yummy;
wire tile_10_4_out_E_noc3_yummy;
wire tile_10_4_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_11_4_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_11_4_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_11_4_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_11_4_out_W_noc1_data;
wire tile_11_4_out_N_noc1_valid;
wire tile_11_4_out_S_noc1_valid;
wire tile_11_4_out_E_noc1_valid;
wire tile_11_4_out_W_noc1_valid;
wire tile_11_4_out_N_noc1_yummy;
wire tile_11_4_out_S_noc1_yummy;
wire tile_11_4_out_E_noc1_yummy;
wire tile_11_4_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_11_4_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_11_4_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_11_4_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_11_4_out_W_noc2_data;
wire tile_11_4_out_N_noc2_valid;
wire tile_11_4_out_S_noc2_valid;
wire tile_11_4_out_E_noc2_valid;
wire tile_11_4_out_W_noc2_valid;
wire tile_11_4_out_N_noc2_yummy;
wire tile_11_4_out_S_noc2_yummy;
wire tile_11_4_out_E_noc2_yummy;
wire tile_11_4_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_11_4_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_11_4_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_11_4_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_11_4_out_W_noc3_data;
wire tile_11_4_out_N_noc3_valid;
wire tile_11_4_out_S_noc3_valid;
wire tile_11_4_out_E_noc3_valid;
wire tile_11_4_out_W_noc3_valid;
wire tile_11_4_out_N_noc3_yummy;
wire tile_11_4_out_S_noc3_yummy;
wire tile_11_4_out_E_noc3_yummy;
wire tile_11_4_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_12_4_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_12_4_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_12_4_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_12_4_out_W_noc1_data;
wire tile_12_4_out_N_noc1_valid;
wire tile_12_4_out_S_noc1_valid;
wire tile_12_4_out_E_noc1_valid;
wire tile_12_4_out_W_noc1_valid;
wire tile_12_4_out_N_noc1_yummy;
wire tile_12_4_out_S_noc1_yummy;
wire tile_12_4_out_E_noc1_yummy;
wire tile_12_4_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_12_4_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_12_4_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_12_4_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_12_4_out_W_noc2_data;
wire tile_12_4_out_N_noc2_valid;
wire tile_12_4_out_S_noc2_valid;
wire tile_12_4_out_E_noc2_valid;
wire tile_12_4_out_W_noc2_valid;
wire tile_12_4_out_N_noc2_yummy;
wire tile_12_4_out_S_noc2_yummy;
wire tile_12_4_out_E_noc2_yummy;
wire tile_12_4_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_12_4_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_12_4_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_12_4_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_12_4_out_W_noc3_data;
wire tile_12_4_out_N_noc3_valid;
wire tile_12_4_out_S_noc3_valid;
wire tile_12_4_out_E_noc3_valid;
wire tile_12_4_out_W_noc3_valid;
wire tile_12_4_out_N_noc3_yummy;
wire tile_12_4_out_S_noc3_yummy;
wire tile_12_4_out_E_noc3_yummy;
wire tile_12_4_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_13_4_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_13_4_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_13_4_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_13_4_out_W_noc1_data;
wire tile_13_4_out_N_noc1_valid;
wire tile_13_4_out_S_noc1_valid;
wire tile_13_4_out_E_noc1_valid;
wire tile_13_4_out_W_noc1_valid;
wire tile_13_4_out_N_noc1_yummy;
wire tile_13_4_out_S_noc1_yummy;
wire tile_13_4_out_E_noc1_yummy;
wire tile_13_4_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_13_4_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_13_4_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_13_4_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_13_4_out_W_noc2_data;
wire tile_13_4_out_N_noc2_valid;
wire tile_13_4_out_S_noc2_valid;
wire tile_13_4_out_E_noc2_valid;
wire tile_13_4_out_W_noc2_valid;
wire tile_13_4_out_N_noc2_yummy;
wire tile_13_4_out_S_noc2_yummy;
wire tile_13_4_out_E_noc2_yummy;
wire tile_13_4_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_13_4_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_13_4_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_13_4_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_13_4_out_W_noc3_data;
wire tile_13_4_out_N_noc3_valid;
wire tile_13_4_out_S_noc3_valid;
wire tile_13_4_out_E_noc3_valid;
wire tile_13_4_out_W_noc3_valid;
wire tile_13_4_out_N_noc3_yummy;
wire tile_13_4_out_S_noc3_yummy;
wire tile_13_4_out_E_noc3_yummy;
wire tile_13_4_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_14_4_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_14_4_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_14_4_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_14_4_out_W_noc1_data;
wire tile_14_4_out_N_noc1_valid;
wire tile_14_4_out_S_noc1_valid;
wire tile_14_4_out_E_noc1_valid;
wire tile_14_4_out_W_noc1_valid;
wire tile_14_4_out_N_noc1_yummy;
wire tile_14_4_out_S_noc1_yummy;
wire tile_14_4_out_E_noc1_yummy;
wire tile_14_4_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_14_4_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_14_4_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_14_4_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_14_4_out_W_noc2_data;
wire tile_14_4_out_N_noc2_valid;
wire tile_14_4_out_S_noc2_valid;
wire tile_14_4_out_E_noc2_valid;
wire tile_14_4_out_W_noc2_valid;
wire tile_14_4_out_N_noc2_yummy;
wire tile_14_4_out_S_noc2_yummy;
wire tile_14_4_out_E_noc2_yummy;
wire tile_14_4_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_14_4_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_14_4_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_14_4_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_14_4_out_W_noc3_data;
wire tile_14_4_out_N_noc3_valid;
wire tile_14_4_out_S_noc3_valid;
wire tile_14_4_out_E_noc3_valid;
wire tile_14_4_out_W_noc3_valid;
wire tile_14_4_out_N_noc3_yummy;
wire tile_14_4_out_S_noc3_yummy;
wire tile_14_4_out_E_noc3_yummy;
wire tile_14_4_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_15_4_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_15_4_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_15_4_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_15_4_out_W_noc1_data;
wire tile_15_4_out_N_noc1_valid;
wire tile_15_4_out_S_noc1_valid;
wire tile_15_4_out_E_noc1_valid;
wire tile_15_4_out_W_noc1_valid;
wire tile_15_4_out_N_noc1_yummy;
wire tile_15_4_out_S_noc1_yummy;
wire tile_15_4_out_E_noc1_yummy;
wire tile_15_4_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_15_4_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_15_4_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_15_4_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_15_4_out_W_noc2_data;
wire tile_15_4_out_N_noc2_valid;
wire tile_15_4_out_S_noc2_valid;
wire tile_15_4_out_E_noc2_valid;
wire tile_15_4_out_W_noc2_valid;
wire tile_15_4_out_N_noc2_yummy;
wire tile_15_4_out_S_noc2_yummy;
wire tile_15_4_out_E_noc2_yummy;
wire tile_15_4_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_15_4_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_15_4_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_15_4_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_15_4_out_W_noc3_data;
wire tile_15_4_out_N_noc3_valid;
wire tile_15_4_out_S_noc3_valid;
wire tile_15_4_out_E_noc3_valid;
wire tile_15_4_out_W_noc3_valid;
wire tile_15_4_out_N_noc3_yummy;
wire tile_15_4_out_S_noc3_yummy;
wire tile_15_4_out_E_noc3_yummy;
wire tile_15_4_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_0_5_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_0_5_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_0_5_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_0_5_out_W_noc1_data;
wire tile_0_5_out_N_noc1_valid;
wire tile_0_5_out_S_noc1_valid;
wire tile_0_5_out_E_noc1_valid;
wire tile_0_5_out_W_noc1_valid;
wire tile_0_5_out_N_noc1_yummy;
wire tile_0_5_out_S_noc1_yummy;
wire tile_0_5_out_E_noc1_yummy;
wire tile_0_5_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_0_5_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_0_5_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_0_5_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_0_5_out_W_noc2_data;
wire tile_0_5_out_N_noc2_valid;
wire tile_0_5_out_S_noc2_valid;
wire tile_0_5_out_E_noc2_valid;
wire tile_0_5_out_W_noc2_valid;
wire tile_0_5_out_N_noc2_yummy;
wire tile_0_5_out_S_noc2_yummy;
wire tile_0_5_out_E_noc2_yummy;
wire tile_0_5_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_0_5_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_0_5_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_0_5_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_0_5_out_W_noc3_data;
wire tile_0_5_out_N_noc3_valid;
wire tile_0_5_out_S_noc3_valid;
wire tile_0_5_out_E_noc3_valid;
wire tile_0_5_out_W_noc3_valid;
wire tile_0_5_out_N_noc3_yummy;
wire tile_0_5_out_S_noc3_yummy;
wire tile_0_5_out_E_noc3_yummy;
wire tile_0_5_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_1_5_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_1_5_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_1_5_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_1_5_out_W_noc1_data;
wire tile_1_5_out_N_noc1_valid;
wire tile_1_5_out_S_noc1_valid;
wire tile_1_5_out_E_noc1_valid;
wire tile_1_5_out_W_noc1_valid;
wire tile_1_5_out_N_noc1_yummy;
wire tile_1_5_out_S_noc1_yummy;
wire tile_1_5_out_E_noc1_yummy;
wire tile_1_5_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_1_5_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_1_5_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_1_5_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_1_5_out_W_noc2_data;
wire tile_1_5_out_N_noc2_valid;
wire tile_1_5_out_S_noc2_valid;
wire tile_1_5_out_E_noc2_valid;
wire tile_1_5_out_W_noc2_valid;
wire tile_1_5_out_N_noc2_yummy;
wire tile_1_5_out_S_noc2_yummy;
wire tile_1_5_out_E_noc2_yummy;
wire tile_1_5_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_1_5_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_1_5_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_1_5_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_1_5_out_W_noc3_data;
wire tile_1_5_out_N_noc3_valid;
wire tile_1_5_out_S_noc3_valid;
wire tile_1_5_out_E_noc3_valid;
wire tile_1_5_out_W_noc3_valid;
wire tile_1_5_out_N_noc3_yummy;
wire tile_1_5_out_S_noc3_yummy;
wire tile_1_5_out_E_noc3_yummy;
wire tile_1_5_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_2_5_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_2_5_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_2_5_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_2_5_out_W_noc1_data;
wire tile_2_5_out_N_noc1_valid;
wire tile_2_5_out_S_noc1_valid;
wire tile_2_5_out_E_noc1_valid;
wire tile_2_5_out_W_noc1_valid;
wire tile_2_5_out_N_noc1_yummy;
wire tile_2_5_out_S_noc1_yummy;
wire tile_2_5_out_E_noc1_yummy;
wire tile_2_5_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_2_5_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_2_5_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_2_5_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_2_5_out_W_noc2_data;
wire tile_2_5_out_N_noc2_valid;
wire tile_2_5_out_S_noc2_valid;
wire tile_2_5_out_E_noc2_valid;
wire tile_2_5_out_W_noc2_valid;
wire tile_2_5_out_N_noc2_yummy;
wire tile_2_5_out_S_noc2_yummy;
wire tile_2_5_out_E_noc2_yummy;
wire tile_2_5_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_2_5_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_2_5_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_2_5_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_2_5_out_W_noc3_data;
wire tile_2_5_out_N_noc3_valid;
wire tile_2_5_out_S_noc3_valid;
wire tile_2_5_out_E_noc3_valid;
wire tile_2_5_out_W_noc3_valid;
wire tile_2_5_out_N_noc3_yummy;
wire tile_2_5_out_S_noc3_yummy;
wire tile_2_5_out_E_noc3_yummy;
wire tile_2_5_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_3_5_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_3_5_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_3_5_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_3_5_out_W_noc1_data;
wire tile_3_5_out_N_noc1_valid;
wire tile_3_5_out_S_noc1_valid;
wire tile_3_5_out_E_noc1_valid;
wire tile_3_5_out_W_noc1_valid;
wire tile_3_5_out_N_noc1_yummy;
wire tile_3_5_out_S_noc1_yummy;
wire tile_3_5_out_E_noc1_yummy;
wire tile_3_5_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_3_5_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_3_5_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_3_5_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_3_5_out_W_noc2_data;
wire tile_3_5_out_N_noc2_valid;
wire tile_3_5_out_S_noc2_valid;
wire tile_3_5_out_E_noc2_valid;
wire tile_3_5_out_W_noc2_valid;
wire tile_3_5_out_N_noc2_yummy;
wire tile_3_5_out_S_noc2_yummy;
wire tile_3_5_out_E_noc2_yummy;
wire tile_3_5_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_3_5_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_3_5_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_3_5_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_3_5_out_W_noc3_data;
wire tile_3_5_out_N_noc3_valid;
wire tile_3_5_out_S_noc3_valid;
wire tile_3_5_out_E_noc3_valid;
wire tile_3_5_out_W_noc3_valid;
wire tile_3_5_out_N_noc3_yummy;
wire tile_3_5_out_S_noc3_yummy;
wire tile_3_5_out_E_noc3_yummy;
wire tile_3_5_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_4_5_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_4_5_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_4_5_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_4_5_out_W_noc1_data;
wire tile_4_5_out_N_noc1_valid;
wire tile_4_5_out_S_noc1_valid;
wire tile_4_5_out_E_noc1_valid;
wire tile_4_5_out_W_noc1_valid;
wire tile_4_5_out_N_noc1_yummy;
wire tile_4_5_out_S_noc1_yummy;
wire tile_4_5_out_E_noc1_yummy;
wire tile_4_5_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_4_5_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_4_5_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_4_5_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_4_5_out_W_noc2_data;
wire tile_4_5_out_N_noc2_valid;
wire tile_4_5_out_S_noc2_valid;
wire tile_4_5_out_E_noc2_valid;
wire tile_4_5_out_W_noc2_valid;
wire tile_4_5_out_N_noc2_yummy;
wire tile_4_5_out_S_noc2_yummy;
wire tile_4_5_out_E_noc2_yummy;
wire tile_4_5_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_4_5_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_4_5_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_4_5_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_4_5_out_W_noc3_data;
wire tile_4_5_out_N_noc3_valid;
wire tile_4_5_out_S_noc3_valid;
wire tile_4_5_out_E_noc3_valid;
wire tile_4_5_out_W_noc3_valid;
wire tile_4_5_out_N_noc3_yummy;
wire tile_4_5_out_S_noc3_yummy;
wire tile_4_5_out_E_noc3_yummy;
wire tile_4_5_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_5_5_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_5_5_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_5_5_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_5_5_out_W_noc1_data;
wire tile_5_5_out_N_noc1_valid;
wire tile_5_5_out_S_noc1_valid;
wire tile_5_5_out_E_noc1_valid;
wire tile_5_5_out_W_noc1_valid;
wire tile_5_5_out_N_noc1_yummy;
wire tile_5_5_out_S_noc1_yummy;
wire tile_5_5_out_E_noc1_yummy;
wire tile_5_5_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_5_5_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_5_5_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_5_5_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_5_5_out_W_noc2_data;
wire tile_5_5_out_N_noc2_valid;
wire tile_5_5_out_S_noc2_valid;
wire tile_5_5_out_E_noc2_valid;
wire tile_5_5_out_W_noc2_valid;
wire tile_5_5_out_N_noc2_yummy;
wire tile_5_5_out_S_noc2_yummy;
wire tile_5_5_out_E_noc2_yummy;
wire tile_5_5_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_5_5_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_5_5_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_5_5_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_5_5_out_W_noc3_data;
wire tile_5_5_out_N_noc3_valid;
wire tile_5_5_out_S_noc3_valid;
wire tile_5_5_out_E_noc3_valid;
wire tile_5_5_out_W_noc3_valid;
wire tile_5_5_out_N_noc3_yummy;
wire tile_5_5_out_S_noc3_yummy;
wire tile_5_5_out_E_noc3_yummy;
wire tile_5_5_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_6_5_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_6_5_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_6_5_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_6_5_out_W_noc1_data;
wire tile_6_5_out_N_noc1_valid;
wire tile_6_5_out_S_noc1_valid;
wire tile_6_5_out_E_noc1_valid;
wire tile_6_5_out_W_noc1_valid;
wire tile_6_5_out_N_noc1_yummy;
wire tile_6_5_out_S_noc1_yummy;
wire tile_6_5_out_E_noc1_yummy;
wire tile_6_5_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_6_5_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_6_5_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_6_5_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_6_5_out_W_noc2_data;
wire tile_6_5_out_N_noc2_valid;
wire tile_6_5_out_S_noc2_valid;
wire tile_6_5_out_E_noc2_valid;
wire tile_6_5_out_W_noc2_valid;
wire tile_6_5_out_N_noc2_yummy;
wire tile_6_5_out_S_noc2_yummy;
wire tile_6_5_out_E_noc2_yummy;
wire tile_6_5_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_6_5_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_6_5_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_6_5_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_6_5_out_W_noc3_data;
wire tile_6_5_out_N_noc3_valid;
wire tile_6_5_out_S_noc3_valid;
wire tile_6_5_out_E_noc3_valid;
wire tile_6_5_out_W_noc3_valid;
wire tile_6_5_out_N_noc3_yummy;
wire tile_6_5_out_S_noc3_yummy;
wire tile_6_5_out_E_noc3_yummy;
wire tile_6_5_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_7_5_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_7_5_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_7_5_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_7_5_out_W_noc1_data;
wire tile_7_5_out_N_noc1_valid;
wire tile_7_5_out_S_noc1_valid;
wire tile_7_5_out_E_noc1_valid;
wire tile_7_5_out_W_noc1_valid;
wire tile_7_5_out_N_noc1_yummy;
wire tile_7_5_out_S_noc1_yummy;
wire tile_7_5_out_E_noc1_yummy;
wire tile_7_5_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_7_5_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_7_5_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_7_5_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_7_5_out_W_noc2_data;
wire tile_7_5_out_N_noc2_valid;
wire tile_7_5_out_S_noc2_valid;
wire tile_7_5_out_E_noc2_valid;
wire tile_7_5_out_W_noc2_valid;
wire tile_7_5_out_N_noc2_yummy;
wire tile_7_5_out_S_noc2_yummy;
wire tile_7_5_out_E_noc2_yummy;
wire tile_7_5_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_7_5_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_7_5_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_7_5_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_7_5_out_W_noc3_data;
wire tile_7_5_out_N_noc3_valid;
wire tile_7_5_out_S_noc3_valid;
wire tile_7_5_out_E_noc3_valid;
wire tile_7_5_out_W_noc3_valid;
wire tile_7_5_out_N_noc3_yummy;
wire tile_7_5_out_S_noc3_yummy;
wire tile_7_5_out_E_noc3_yummy;
wire tile_7_5_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_8_5_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_8_5_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_8_5_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_8_5_out_W_noc1_data;
wire tile_8_5_out_N_noc1_valid;
wire tile_8_5_out_S_noc1_valid;
wire tile_8_5_out_E_noc1_valid;
wire tile_8_5_out_W_noc1_valid;
wire tile_8_5_out_N_noc1_yummy;
wire tile_8_5_out_S_noc1_yummy;
wire tile_8_5_out_E_noc1_yummy;
wire tile_8_5_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_8_5_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_8_5_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_8_5_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_8_5_out_W_noc2_data;
wire tile_8_5_out_N_noc2_valid;
wire tile_8_5_out_S_noc2_valid;
wire tile_8_5_out_E_noc2_valid;
wire tile_8_5_out_W_noc2_valid;
wire tile_8_5_out_N_noc2_yummy;
wire tile_8_5_out_S_noc2_yummy;
wire tile_8_5_out_E_noc2_yummy;
wire tile_8_5_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_8_5_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_8_5_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_8_5_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_8_5_out_W_noc3_data;
wire tile_8_5_out_N_noc3_valid;
wire tile_8_5_out_S_noc3_valid;
wire tile_8_5_out_E_noc3_valid;
wire tile_8_5_out_W_noc3_valid;
wire tile_8_5_out_N_noc3_yummy;
wire tile_8_5_out_S_noc3_yummy;
wire tile_8_5_out_E_noc3_yummy;
wire tile_8_5_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_9_5_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_9_5_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_9_5_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_9_5_out_W_noc1_data;
wire tile_9_5_out_N_noc1_valid;
wire tile_9_5_out_S_noc1_valid;
wire tile_9_5_out_E_noc1_valid;
wire tile_9_5_out_W_noc1_valid;
wire tile_9_5_out_N_noc1_yummy;
wire tile_9_5_out_S_noc1_yummy;
wire tile_9_5_out_E_noc1_yummy;
wire tile_9_5_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_9_5_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_9_5_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_9_5_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_9_5_out_W_noc2_data;
wire tile_9_5_out_N_noc2_valid;
wire tile_9_5_out_S_noc2_valid;
wire tile_9_5_out_E_noc2_valid;
wire tile_9_5_out_W_noc2_valid;
wire tile_9_5_out_N_noc2_yummy;
wire tile_9_5_out_S_noc2_yummy;
wire tile_9_5_out_E_noc2_yummy;
wire tile_9_5_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_9_5_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_9_5_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_9_5_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_9_5_out_W_noc3_data;
wire tile_9_5_out_N_noc3_valid;
wire tile_9_5_out_S_noc3_valid;
wire tile_9_5_out_E_noc3_valid;
wire tile_9_5_out_W_noc3_valid;
wire tile_9_5_out_N_noc3_yummy;
wire tile_9_5_out_S_noc3_yummy;
wire tile_9_5_out_E_noc3_yummy;
wire tile_9_5_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_10_5_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_10_5_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_10_5_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_10_5_out_W_noc1_data;
wire tile_10_5_out_N_noc1_valid;
wire tile_10_5_out_S_noc1_valid;
wire tile_10_5_out_E_noc1_valid;
wire tile_10_5_out_W_noc1_valid;
wire tile_10_5_out_N_noc1_yummy;
wire tile_10_5_out_S_noc1_yummy;
wire tile_10_5_out_E_noc1_yummy;
wire tile_10_5_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_10_5_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_10_5_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_10_5_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_10_5_out_W_noc2_data;
wire tile_10_5_out_N_noc2_valid;
wire tile_10_5_out_S_noc2_valid;
wire tile_10_5_out_E_noc2_valid;
wire tile_10_5_out_W_noc2_valid;
wire tile_10_5_out_N_noc2_yummy;
wire tile_10_5_out_S_noc2_yummy;
wire tile_10_5_out_E_noc2_yummy;
wire tile_10_5_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_10_5_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_10_5_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_10_5_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_10_5_out_W_noc3_data;
wire tile_10_5_out_N_noc3_valid;
wire tile_10_5_out_S_noc3_valid;
wire tile_10_5_out_E_noc3_valid;
wire tile_10_5_out_W_noc3_valid;
wire tile_10_5_out_N_noc3_yummy;
wire tile_10_5_out_S_noc3_yummy;
wire tile_10_5_out_E_noc3_yummy;
wire tile_10_5_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_11_5_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_11_5_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_11_5_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_11_5_out_W_noc1_data;
wire tile_11_5_out_N_noc1_valid;
wire tile_11_5_out_S_noc1_valid;
wire tile_11_5_out_E_noc1_valid;
wire tile_11_5_out_W_noc1_valid;
wire tile_11_5_out_N_noc1_yummy;
wire tile_11_5_out_S_noc1_yummy;
wire tile_11_5_out_E_noc1_yummy;
wire tile_11_5_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_11_5_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_11_5_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_11_5_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_11_5_out_W_noc2_data;
wire tile_11_5_out_N_noc2_valid;
wire tile_11_5_out_S_noc2_valid;
wire tile_11_5_out_E_noc2_valid;
wire tile_11_5_out_W_noc2_valid;
wire tile_11_5_out_N_noc2_yummy;
wire tile_11_5_out_S_noc2_yummy;
wire tile_11_5_out_E_noc2_yummy;
wire tile_11_5_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_11_5_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_11_5_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_11_5_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_11_5_out_W_noc3_data;
wire tile_11_5_out_N_noc3_valid;
wire tile_11_5_out_S_noc3_valid;
wire tile_11_5_out_E_noc3_valid;
wire tile_11_5_out_W_noc3_valid;
wire tile_11_5_out_N_noc3_yummy;
wire tile_11_5_out_S_noc3_yummy;
wire tile_11_5_out_E_noc3_yummy;
wire tile_11_5_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_12_5_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_12_5_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_12_5_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_12_5_out_W_noc1_data;
wire tile_12_5_out_N_noc1_valid;
wire tile_12_5_out_S_noc1_valid;
wire tile_12_5_out_E_noc1_valid;
wire tile_12_5_out_W_noc1_valid;
wire tile_12_5_out_N_noc1_yummy;
wire tile_12_5_out_S_noc1_yummy;
wire tile_12_5_out_E_noc1_yummy;
wire tile_12_5_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_12_5_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_12_5_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_12_5_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_12_5_out_W_noc2_data;
wire tile_12_5_out_N_noc2_valid;
wire tile_12_5_out_S_noc2_valid;
wire tile_12_5_out_E_noc2_valid;
wire tile_12_5_out_W_noc2_valid;
wire tile_12_5_out_N_noc2_yummy;
wire tile_12_5_out_S_noc2_yummy;
wire tile_12_5_out_E_noc2_yummy;
wire tile_12_5_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_12_5_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_12_5_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_12_5_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_12_5_out_W_noc3_data;
wire tile_12_5_out_N_noc3_valid;
wire tile_12_5_out_S_noc3_valid;
wire tile_12_5_out_E_noc3_valid;
wire tile_12_5_out_W_noc3_valid;
wire tile_12_5_out_N_noc3_yummy;
wire tile_12_5_out_S_noc3_yummy;
wire tile_12_5_out_E_noc3_yummy;
wire tile_12_5_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_13_5_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_13_5_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_13_5_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_13_5_out_W_noc1_data;
wire tile_13_5_out_N_noc1_valid;
wire tile_13_5_out_S_noc1_valid;
wire tile_13_5_out_E_noc1_valid;
wire tile_13_5_out_W_noc1_valid;
wire tile_13_5_out_N_noc1_yummy;
wire tile_13_5_out_S_noc1_yummy;
wire tile_13_5_out_E_noc1_yummy;
wire tile_13_5_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_13_5_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_13_5_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_13_5_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_13_5_out_W_noc2_data;
wire tile_13_5_out_N_noc2_valid;
wire tile_13_5_out_S_noc2_valid;
wire tile_13_5_out_E_noc2_valid;
wire tile_13_5_out_W_noc2_valid;
wire tile_13_5_out_N_noc2_yummy;
wire tile_13_5_out_S_noc2_yummy;
wire tile_13_5_out_E_noc2_yummy;
wire tile_13_5_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_13_5_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_13_5_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_13_5_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_13_5_out_W_noc3_data;
wire tile_13_5_out_N_noc3_valid;
wire tile_13_5_out_S_noc3_valid;
wire tile_13_5_out_E_noc3_valid;
wire tile_13_5_out_W_noc3_valid;
wire tile_13_5_out_N_noc3_yummy;
wire tile_13_5_out_S_noc3_yummy;
wire tile_13_5_out_E_noc3_yummy;
wire tile_13_5_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_14_5_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_14_5_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_14_5_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_14_5_out_W_noc1_data;
wire tile_14_5_out_N_noc1_valid;
wire tile_14_5_out_S_noc1_valid;
wire tile_14_5_out_E_noc1_valid;
wire tile_14_5_out_W_noc1_valid;
wire tile_14_5_out_N_noc1_yummy;
wire tile_14_5_out_S_noc1_yummy;
wire tile_14_5_out_E_noc1_yummy;
wire tile_14_5_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_14_5_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_14_5_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_14_5_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_14_5_out_W_noc2_data;
wire tile_14_5_out_N_noc2_valid;
wire tile_14_5_out_S_noc2_valid;
wire tile_14_5_out_E_noc2_valid;
wire tile_14_5_out_W_noc2_valid;
wire tile_14_5_out_N_noc2_yummy;
wire tile_14_5_out_S_noc2_yummy;
wire tile_14_5_out_E_noc2_yummy;
wire tile_14_5_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_14_5_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_14_5_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_14_5_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_14_5_out_W_noc3_data;
wire tile_14_5_out_N_noc3_valid;
wire tile_14_5_out_S_noc3_valid;
wire tile_14_5_out_E_noc3_valid;
wire tile_14_5_out_W_noc3_valid;
wire tile_14_5_out_N_noc3_yummy;
wire tile_14_5_out_S_noc3_yummy;
wire tile_14_5_out_E_noc3_yummy;
wire tile_14_5_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_15_5_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_15_5_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_15_5_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_15_5_out_W_noc1_data;
wire tile_15_5_out_N_noc1_valid;
wire tile_15_5_out_S_noc1_valid;
wire tile_15_5_out_E_noc1_valid;
wire tile_15_5_out_W_noc1_valid;
wire tile_15_5_out_N_noc1_yummy;
wire tile_15_5_out_S_noc1_yummy;
wire tile_15_5_out_E_noc1_yummy;
wire tile_15_5_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_15_5_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_15_5_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_15_5_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_15_5_out_W_noc2_data;
wire tile_15_5_out_N_noc2_valid;
wire tile_15_5_out_S_noc2_valid;
wire tile_15_5_out_E_noc2_valid;
wire tile_15_5_out_W_noc2_valid;
wire tile_15_5_out_N_noc2_yummy;
wire tile_15_5_out_S_noc2_yummy;
wire tile_15_5_out_E_noc2_yummy;
wire tile_15_5_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_15_5_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_15_5_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_15_5_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_15_5_out_W_noc3_data;
wire tile_15_5_out_N_noc3_valid;
wire tile_15_5_out_S_noc3_valid;
wire tile_15_5_out_E_noc3_valid;
wire tile_15_5_out_W_noc3_valid;
wire tile_15_5_out_N_noc3_yummy;
wire tile_15_5_out_S_noc3_yummy;
wire tile_15_5_out_E_noc3_yummy;
wire tile_15_5_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_0_6_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_0_6_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_0_6_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_0_6_out_W_noc1_data;
wire tile_0_6_out_N_noc1_valid;
wire tile_0_6_out_S_noc1_valid;
wire tile_0_6_out_E_noc1_valid;
wire tile_0_6_out_W_noc1_valid;
wire tile_0_6_out_N_noc1_yummy;
wire tile_0_6_out_S_noc1_yummy;
wire tile_0_6_out_E_noc1_yummy;
wire tile_0_6_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_0_6_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_0_6_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_0_6_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_0_6_out_W_noc2_data;
wire tile_0_6_out_N_noc2_valid;
wire tile_0_6_out_S_noc2_valid;
wire tile_0_6_out_E_noc2_valid;
wire tile_0_6_out_W_noc2_valid;
wire tile_0_6_out_N_noc2_yummy;
wire tile_0_6_out_S_noc2_yummy;
wire tile_0_6_out_E_noc2_yummy;
wire tile_0_6_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_0_6_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_0_6_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_0_6_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_0_6_out_W_noc3_data;
wire tile_0_6_out_N_noc3_valid;
wire tile_0_6_out_S_noc3_valid;
wire tile_0_6_out_E_noc3_valid;
wire tile_0_6_out_W_noc3_valid;
wire tile_0_6_out_N_noc3_yummy;
wire tile_0_6_out_S_noc3_yummy;
wire tile_0_6_out_E_noc3_yummy;
wire tile_0_6_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_1_6_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_1_6_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_1_6_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_1_6_out_W_noc1_data;
wire tile_1_6_out_N_noc1_valid;
wire tile_1_6_out_S_noc1_valid;
wire tile_1_6_out_E_noc1_valid;
wire tile_1_6_out_W_noc1_valid;
wire tile_1_6_out_N_noc1_yummy;
wire tile_1_6_out_S_noc1_yummy;
wire tile_1_6_out_E_noc1_yummy;
wire tile_1_6_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_1_6_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_1_6_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_1_6_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_1_6_out_W_noc2_data;
wire tile_1_6_out_N_noc2_valid;
wire tile_1_6_out_S_noc2_valid;
wire tile_1_6_out_E_noc2_valid;
wire tile_1_6_out_W_noc2_valid;
wire tile_1_6_out_N_noc2_yummy;
wire tile_1_6_out_S_noc2_yummy;
wire tile_1_6_out_E_noc2_yummy;
wire tile_1_6_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_1_6_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_1_6_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_1_6_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_1_6_out_W_noc3_data;
wire tile_1_6_out_N_noc3_valid;
wire tile_1_6_out_S_noc3_valid;
wire tile_1_6_out_E_noc3_valid;
wire tile_1_6_out_W_noc3_valid;
wire tile_1_6_out_N_noc3_yummy;
wire tile_1_6_out_S_noc3_yummy;
wire tile_1_6_out_E_noc3_yummy;
wire tile_1_6_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_2_6_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_2_6_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_2_6_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_2_6_out_W_noc1_data;
wire tile_2_6_out_N_noc1_valid;
wire tile_2_6_out_S_noc1_valid;
wire tile_2_6_out_E_noc1_valid;
wire tile_2_6_out_W_noc1_valid;
wire tile_2_6_out_N_noc1_yummy;
wire tile_2_6_out_S_noc1_yummy;
wire tile_2_6_out_E_noc1_yummy;
wire tile_2_6_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_2_6_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_2_6_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_2_6_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_2_6_out_W_noc2_data;
wire tile_2_6_out_N_noc2_valid;
wire tile_2_6_out_S_noc2_valid;
wire tile_2_6_out_E_noc2_valid;
wire tile_2_6_out_W_noc2_valid;
wire tile_2_6_out_N_noc2_yummy;
wire tile_2_6_out_S_noc2_yummy;
wire tile_2_6_out_E_noc2_yummy;
wire tile_2_6_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_2_6_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_2_6_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_2_6_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_2_6_out_W_noc3_data;
wire tile_2_6_out_N_noc3_valid;
wire tile_2_6_out_S_noc3_valid;
wire tile_2_6_out_E_noc3_valid;
wire tile_2_6_out_W_noc3_valid;
wire tile_2_6_out_N_noc3_yummy;
wire tile_2_6_out_S_noc3_yummy;
wire tile_2_6_out_E_noc3_yummy;
wire tile_2_6_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_3_6_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_3_6_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_3_6_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_3_6_out_W_noc1_data;
wire tile_3_6_out_N_noc1_valid;
wire tile_3_6_out_S_noc1_valid;
wire tile_3_6_out_E_noc1_valid;
wire tile_3_6_out_W_noc1_valid;
wire tile_3_6_out_N_noc1_yummy;
wire tile_3_6_out_S_noc1_yummy;
wire tile_3_6_out_E_noc1_yummy;
wire tile_3_6_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_3_6_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_3_6_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_3_6_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_3_6_out_W_noc2_data;
wire tile_3_6_out_N_noc2_valid;
wire tile_3_6_out_S_noc2_valid;
wire tile_3_6_out_E_noc2_valid;
wire tile_3_6_out_W_noc2_valid;
wire tile_3_6_out_N_noc2_yummy;
wire tile_3_6_out_S_noc2_yummy;
wire tile_3_6_out_E_noc2_yummy;
wire tile_3_6_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_3_6_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_3_6_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_3_6_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_3_6_out_W_noc3_data;
wire tile_3_6_out_N_noc3_valid;
wire tile_3_6_out_S_noc3_valid;
wire tile_3_6_out_E_noc3_valid;
wire tile_3_6_out_W_noc3_valid;
wire tile_3_6_out_N_noc3_yummy;
wire tile_3_6_out_S_noc3_yummy;
wire tile_3_6_out_E_noc3_yummy;
wire tile_3_6_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_4_6_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_4_6_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_4_6_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_4_6_out_W_noc1_data;
wire tile_4_6_out_N_noc1_valid;
wire tile_4_6_out_S_noc1_valid;
wire tile_4_6_out_E_noc1_valid;
wire tile_4_6_out_W_noc1_valid;
wire tile_4_6_out_N_noc1_yummy;
wire tile_4_6_out_S_noc1_yummy;
wire tile_4_6_out_E_noc1_yummy;
wire tile_4_6_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_4_6_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_4_6_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_4_6_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_4_6_out_W_noc2_data;
wire tile_4_6_out_N_noc2_valid;
wire tile_4_6_out_S_noc2_valid;
wire tile_4_6_out_E_noc2_valid;
wire tile_4_6_out_W_noc2_valid;
wire tile_4_6_out_N_noc2_yummy;
wire tile_4_6_out_S_noc2_yummy;
wire tile_4_6_out_E_noc2_yummy;
wire tile_4_6_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_4_6_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_4_6_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_4_6_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_4_6_out_W_noc3_data;
wire tile_4_6_out_N_noc3_valid;
wire tile_4_6_out_S_noc3_valid;
wire tile_4_6_out_E_noc3_valid;
wire tile_4_6_out_W_noc3_valid;
wire tile_4_6_out_N_noc3_yummy;
wire tile_4_6_out_S_noc3_yummy;
wire tile_4_6_out_E_noc3_yummy;
wire tile_4_6_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_5_6_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_5_6_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_5_6_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_5_6_out_W_noc1_data;
wire tile_5_6_out_N_noc1_valid;
wire tile_5_6_out_S_noc1_valid;
wire tile_5_6_out_E_noc1_valid;
wire tile_5_6_out_W_noc1_valid;
wire tile_5_6_out_N_noc1_yummy;
wire tile_5_6_out_S_noc1_yummy;
wire tile_5_6_out_E_noc1_yummy;
wire tile_5_6_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_5_6_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_5_6_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_5_6_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_5_6_out_W_noc2_data;
wire tile_5_6_out_N_noc2_valid;
wire tile_5_6_out_S_noc2_valid;
wire tile_5_6_out_E_noc2_valid;
wire tile_5_6_out_W_noc2_valid;
wire tile_5_6_out_N_noc2_yummy;
wire tile_5_6_out_S_noc2_yummy;
wire tile_5_6_out_E_noc2_yummy;
wire tile_5_6_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_5_6_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_5_6_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_5_6_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_5_6_out_W_noc3_data;
wire tile_5_6_out_N_noc3_valid;
wire tile_5_6_out_S_noc3_valid;
wire tile_5_6_out_E_noc3_valid;
wire tile_5_6_out_W_noc3_valid;
wire tile_5_6_out_N_noc3_yummy;
wire tile_5_6_out_S_noc3_yummy;
wire tile_5_6_out_E_noc3_yummy;
wire tile_5_6_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_6_6_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_6_6_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_6_6_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_6_6_out_W_noc1_data;
wire tile_6_6_out_N_noc1_valid;
wire tile_6_6_out_S_noc1_valid;
wire tile_6_6_out_E_noc1_valid;
wire tile_6_6_out_W_noc1_valid;
wire tile_6_6_out_N_noc1_yummy;
wire tile_6_6_out_S_noc1_yummy;
wire tile_6_6_out_E_noc1_yummy;
wire tile_6_6_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_6_6_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_6_6_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_6_6_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_6_6_out_W_noc2_data;
wire tile_6_6_out_N_noc2_valid;
wire tile_6_6_out_S_noc2_valid;
wire tile_6_6_out_E_noc2_valid;
wire tile_6_6_out_W_noc2_valid;
wire tile_6_6_out_N_noc2_yummy;
wire tile_6_6_out_S_noc2_yummy;
wire tile_6_6_out_E_noc2_yummy;
wire tile_6_6_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_6_6_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_6_6_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_6_6_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_6_6_out_W_noc3_data;
wire tile_6_6_out_N_noc3_valid;
wire tile_6_6_out_S_noc3_valid;
wire tile_6_6_out_E_noc3_valid;
wire tile_6_6_out_W_noc3_valid;
wire tile_6_6_out_N_noc3_yummy;
wire tile_6_6_out_S_noc3_yummy;
wire tile_6_6_out_E_noc3_yummy;
wire tile_6_6_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_7_6_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_7_6_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_7_6_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_7_6_out_W_noc1_data;
wire tile_7_6_out_N_noc1_valid;
wire tile_7_6_out_S_noc1_valid;
wire tile_7_6_out_E_noc1_valid;
wire tile_7_6_out_W_noc1_valid;
wire tile_7_6_out_N_noc1_yummy;
wire tile_7_6_out_S_noc1_yummy;
wire tile_7_6_out_E_noc1_yummy;
wire tile_7_6_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_7_6_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_7_6_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_7_6_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_7_6_out_W_noc2_data;
wire tile_7_6_out_N_noc2_valid;
wire tile_7_6_out_S_noc2_valid;
wire tile_7_6_out_E_noc2_valid;
wire tile_7_6_out_W_noc2_valid;
wire tile_7_6_out_N_noc2_yummy;
wire tile_7_6_out_S_noc2_yummy;
wire tile_7_6_out_E_noc2_yummy;
wire tile_7_6_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_7_6_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_7_6_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_7_6_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_7_6_out_W_noc3_data;
wire tile_7_6_out_N_noc3_valid;
wire tile_7_6_out_S_noc3_valid;
wire tile_7_6_out_E_noc3_valid;
wire tile_7_6_out_W_noc3_valid;
wire tile_7_6_out_N_noc3_yummy;
wire tile_7_6_out_S_noc3_yummy;
wire tile_7_6_out_E_noc3_yummy;
wire tile_7_6_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_8_6_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_8_6_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_8_6_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_8_6_out_W_noc1_data;
wire tile_8_6_out_N_noc1_valid;
wire tile_8_6_out_S_noc1_valid;
wire tile_8_6_out_E_noc1_valid;
wire tile_8_6_out_W_noc1_valid;
wire tile_8_6_out_N_noc1_yummy;
wire tile_8_6_out_S_noc1_yummy;
wire tile_8_6_out_E_noc1_yummy;
wire tile_8_6_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_8_6_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_8_6_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_8_6_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_8_6_out_W_noc2_data;
wire tile_8_6_out_N_noc2_valid;
wire tile_8_6_out_S_noc2_valid;
wire tile_8_6_out_E_noc2_valid;
wire tile_8_6_out_W_noc2_valid;
wire tile_8_6_out_N_noc2_yummy;
wire tile_8_6_out_S_noc2_yummy;
wire tile_8_6_out_E_noc2_yummy;
wire tile_8_6_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_8_6_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_8_6_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_8_6_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_8_6_out_W_noc3_data;
wire tile_8_6_out_N_noc3_valid;
wire tile_8_6_out_S_noc3_valid;
wire tile_8_6_out_E_noc3_valid;
wire tile_8_6_out_W_noc3_valid;
wire tile_8_6_out_N_noc3_yummy;
wire tile_8_6_out_S_noc3_yummy;
wire tile_8_6_out_E_noc3_yummy;
wire tile_8_6_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_9_6_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_9_6_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_9_6_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_9_6_out_W_noc1_data;
wire tile_9_6_out_N_noc1_valid;
wire tile_9_6_out_S_noc1_valid;
wire tile_9_6_out_E_noc1_valid;
wire tile_9_6_out_W_noc1_valid;
wire tile_9_6_out_N_noc1_yummy;
wire tile_9_6_out_S_noc1_yummy;
wire tile_9_6_out_E_noc1_yummy;
wire tile_9_6_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_9_6_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_9_6_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_9_6_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_9_6_out_W_noc2_data;
wire tile_9_6_out_N_noc2_valid;
wire tile_9_6_out_S_noc2_valid;
wire tile_9_6_out_E_noc2_valid;
wire tile_9_6_out_W_noc2_valid;
wire tile_9_6_out_N_noc2_yummy;
wire tile_9_6_out_S_noc2_yummy;
wire tile_9_6_out_E_noc2_yummy;
wire tile_9_6_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_9_6_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_9_6_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_9_6_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_9_6_out_W_noc3_data;
wire tile_9_6_out_N_noc3_valid;
wire tile_9_6_out_S_noc3_valid;
wire tile_9_6_out_E_noc3_valid;
wire tile_9_6_out_W_noc3_valid;
wire tile_9_6_out_N_noc3_yummy;
wire tile_9_6_out_S_noc3_yummy;
wire tile_9_6_out_E_noc3_yummy;
wire tile_9_6_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_10_6_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_10_6_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_10_6_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_10_6_out_W_noc1_data;
wire tile_10_6_out_N_noc1_valid;
wire tile_10_6_out_S_noc1_valid;
wire tile_10_6_out_E_noc1_valid;
wire tile_10_6_out_W_noc1_valid;
wire tile_10_6_out_N_noc1_yummy;
wire tile_10_6_out_S_noc1_yummy;
wire tile_10_6_out_E_noc1_yummy;
wire tile_10_6_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_10_6_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_10_6_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_10_6_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_10_6_out_W_noc2_data;
wire tile_10_6_out_N_noc2_valid;
wire tile_10_6_out_S_noc2_valid;
wire tile_10_6_out_E_noc2_valid;
wire tile_10_6_out_W_noc2_valid;
wire tile_10_6_out_N_noc2_yummy;
wire tile_10_6_out_S_noc2_yummy;
wire tile_10_6_out_E_noc2_yummy;
wire tile_10_6_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_10_6_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_10_6_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_10_6_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_10_6_out_W_noc3_data;
wire tile_10_6_out_N_noc3_valid;
wire tile_10_6_out_S_noc3_valid;
wire tile_10_6_out_E_noc3_valid;
wire tile_10_6_out_W_noc3_valid;
wire tile_10_6_out_N_noc3_yummy;
wire tile_10_6_out_S_noc3_yummy;
wire tile_10_6_out_E_noc3_yummy;
wire tile_10_6_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_11_6_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_11_6_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_11_6_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_11_6_out_W_noc1_data;
wire tile_11_6_out_N_noc1_valid;
wire tile_11_6_out_S_noc1_valid;
wire tile_11_6_out_E_noc1_valid;
wire tile_11_6_out_W_noc1_valid;
wire tile_11_6_out_N_noc1_yummy;
wire tile_11_6_out_S_noc1_yummy;
wire tile_11_6_out_E_noc1_yummy;
wire tile_11_6_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_11_6_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_11_6_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_11_6_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_11_6_out_W_noc2_data;
wire tile_11_6_out_N_noc2_valid;
wire tile_11_6_out_S_noc2_valid;
wire tile_11_6_out_E_noc2_valid;
wire tile_11_6_out_W_noc2_valid;
wire tile_11_6_out_N_noc2_yummy;
wire tile_11_6_out_S_noc2_yummy;
wire tile_11_6_out_E_noc2_yummy;
wire tile_11_6_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_11_6_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_11_6_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_11_6_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_11_6_out_W_noc3_data;
wire tile_11_6_out_N_noc3_valid;
wire tile_11_6_out_S_noc3_valid;
wire tile_11_6_out_E_noc3_valid;
wire tile_11_6_out_W_noc3_valid;
wire tile_11_6_out_N_noc3_yummy;
wire tile_11_6_out_S_noc3_yummy;
wire tile_11_6_out_E_noc3_yummy;
wire tile_11_6_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_12_6_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_12_6_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_12_6_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_12_6_out_W_noc1_data;
wire tile_12_6_out_N_noc1_valid;
wire tile_12_6_out_S_noc1_valid;
wire tile_12_6_out_E_noc1_valid;
wire tile_12_6_out_W_noc1_valid;
wire tile_12_6_out_N_noc1_yummy;
wire tile_12_6_out_S_noc1_yummy;
wire tile_12_6_out_E_noc1_yummy;
wire tile_12_6_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_12_6_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_12_6_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_12_6_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_12_6_out_W_noc2_data;
wire tile_12_6_out_N_noc2_valid;
wire tile_12_6_out_S_noc2_valid;
wire tile_12_6_out_E_noc2_valid;
wire tile_12_6_out_W_noc2_valid;
wire tile_12_6_out_N_noc2_yummy;
wire tile_12_6_out_S_noc2_yummy;
wire tile_12_6_out_E_noc2_yummy;
wire tile_12_6_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_12_6_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_12_6_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_12_6_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_12_6_out_W_noc3_data;
wire tile_12_6_out_N_noc3_valid;
wire tile_12_6_out_S_noc3_valid;
wire tile_12_6_out_E_noc3_valid;
wire tile_12_6_out_W_noc3_valid;
wire tile_12_6_out_N_noc3_yummy;
wire tile_12_6_out_S_noc3_yummy;
wire tile_12_6_out_E_noc3_yummy;
wire tile_12_6_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_13_6_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_13_6_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_13_6_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_13_6_out_W_noc1_data;
wire tile_13_6_out_N_noc1_valid;
wire tile_13_6_out_S_noc1_valid;
wire tile_13_6_out_E_noc1_valid;
wire tile_13_6_out_W_noc1_valid;
wire tile_13_6_out_N_noc1_yummy;
wire tile_13_6_out_S_noc1_yummy;
wire tile_13_6_out_E_noc1_yummy;
wire tile_13_6_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_13_6_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_13_6_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_13_6_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_13_6_out_W_noc2_data;
wire tile_13_6_out_N_noc2_valid;
wire tile_13_6_out_S_noc2_valid;
wire tile_13_6_out_E_noc2_valid;
wire tile_13_6_out_W_noc2_valid;
wire tile_13_6_out_N_noc2_yummy;
wire tile_13_6_out_S_noc2_yummy;
wire tile_13_6_out_E_noc2_yummy;
wire tile_13_6_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_13_6_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_13_6_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_13_6_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_13_6_out_W_noc3_data;
wire tile_13_6_out_N_noc3_valid;
wire tile_13_6_out_S_noc3_valid;
wire tile_13_6_out_E_noc3_valid;
wire tile_13_6_out_W_noc3_valid;
wire tile_13_6_out_N_noc3_yummy;
wire tile_13_6_out_S_noc3_yummy;
wire tile_13_6_out_E_noc3_yummy;
wire tile_13_6_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_14_6_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_14_6_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_14_6_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_14_6_out_W_noc1_data;
wire tile_14_6_out_N_noc1_valid;
wire tile_14_6_out_S_noc1_valid;
wire tile_14_6_out_E_noc1_valid;
wire tile_14_6_out_W_noc1_valid;
wire tile_14_6_out_N_noc1_yummy;
wire tile_14_6_out_S_noc1_yummy;
wire tile_14_6_out_E_noc1_yummy;
wire tile_14_6_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_14_6_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_14_6_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_14_6_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_14_6_out_W_noc2_data;
wire tile_14_6_out_N_noc2_valid;
wire tile_14_6_out_S_noc2_valid;
wire tile_14_6_out_E_noc2_valid;
wire tile_14_6_out_W_noc2_valid;
wire tile_14_6_out_N_noc2_yummy;
wire tile_14_6_out_S_noc2_yummy;
wire tile_14_6_out_E_noc2_yummy;
wire tile_14_6_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_14_6_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_14_6_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_14_6_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_14_6_out_W_noc3_data;
wire tile_14_6_out_N_noc3_valid;
wire tile_14_6_out_S_noc3_valid;
wire tile_14_6_out_E_noc3_valid;
wire tile_14_6_out_W_noc3_valid;
wire tile_14_6_out_N_noc3_yummy;
wire tile_14_6_out_S_noc3_yummy;
wire tile_14_6_out_E_noc3_yummy;
wire tile_14_6_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_15_6_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_15_6_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_15_6_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_15_6_out_W_noc1_data;
wire tile_15_6_out_N_noc1_valid;
wire tile_15_6_out_S_noc1_valid;
wire tile_15_6_out_E_noc1_valid;
wire tile_15_6_out_W_noc1_valid;
wire tile_15_6_out_N_noc1_yummy;
wire tile_15_6_out_S_noc1_yummy;
wire tile_15_6_out_E_noc1_yummy;
wire tile_15_6_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_15_6_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_15_6_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_15_6_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_15_6_out_W_noc2_data;
wire tile_15_6_out_N_noc2_valid;
wire tile_15_6_out_S_noc2_valid;
wire tile_15_6_out_E_noc2_valid;
wire tile_15_6_out_W_noc2_valid;
wire tile_15_6_out_N_noc2_yummy;
wire tile_15_6_out_S_noc2_yummy;
wire tile_15_6_out_E_noc2_yummy;
wire tile_15_6_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_15_6_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_15_6_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_15_6_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_15_6_out_W_noc3_data;
wire tile_15_6_out_N_noc3_valid;
wire tile_15_6_out_S_noc3_valid;
wire tile_15_6_out_E_noc3_valid;
wire tile_15_6_out_W_noc3_valid;
wire tile_15_6_out_N_noc3_yummy;
wire tile_15_6_out_S_noc3_yummy;
wire tile_15_6_out_E_noc3_yummy;
wire tile_15_6_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_0_7_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_0_7_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_0_7_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_0_7_out_W_noc1_data;
wire tile_0_7_out_N_noc1_valid;
wire tile_0_7_out_S_noc1_valid;
wire tile_0_7_out_E_noc1_valid;
wire tile_0_7_out_W_noc1_valid;
wire tile_0_7_out_N_noc1_yummy;
wire tile_0_7_out_S_noc1_yummy;
wire tile_0_7_out_E_noc1_yummy;
wire tile_0_7_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_0_7_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_0_7_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_0_7_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_0_7_out_W_noc2_data;
wire tile_0_7_out_N_noc2_valid;
wire tile_0_7_out_S_noc2_valid;
wire tile_0_7_out_E_noc2_valid;
wire tile_0_7_out_W_noc2_valid;
wire tile_0_7_out_N_noc2_yummy;
wire tile_0_7_out_S_noc2_yummy;
wire tile_0_7_out_E_noc2_yummy;
wire tile_0_7_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_0_7_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_0_7_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_0_7_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_0_7_out_W_noc3_data;
wire tile_0_7_out_N_noc3_valid;
wire tile_0_7_out_S_noc3_valid;
wire tile_0_7_out_E_noc3_valid;
wire tile_0_7_out_W_noc3_valid;
wire tile_0_7_out_N_noc3_yummy;
wire tile_0_7_out_S_noc3_yummy;
wire tile_0_7_out_E_noc3_yummy;
wire tile_0_7_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_1_7_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_1_7_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_1_7_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_1_7_out_W_noc1_data;
wire tile_1_7_out_N_noc1_valid;
wire tile_1_7_out_S_noc1_valid;
wire tile_1_7_out_E_noc1_valid;
wire tile_1_7_out_W_noc1_valid;
wire tile_1_7_out_N_noc1_yummy;
wire tile_1_7_out_S_noc1_yummy;
wire tile_1_7_out_E_noc1_yummy;
wire tile_1_7_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_1_7_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_1_7_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_1_7_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_1_7_out_W_noc2_data;
wire tile_1_7_out_N_noc2_valid;
wire tile_1_7_out_S_noc2_valid;
wire tile_1_7_out_E_noc2_valid;
wire tile_1_7_out_W_noc2_valid;
wire tile_1_7_out_N_noc2_yummy;
wire tile_1_7_out_S_noc2_yummy;
wire tile_1_7_out_E_noc2_yummy;
wire tile_1_7_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_1_7_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_1_7_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_1_7_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_1_7_out_W_noc3_data;
wire tile_1_7_out_N_noc3_valid;
wire tile_1_7_out_S_noc3_valid;
wire tile_1_7_out_E_noc3_valid;
wire tile_1_7_out_W_noc3_valid;
wire tile_1_7_out_N_noc3_yummy;
wire tile_1_7_out_S_noc3_yummy;
wire tile_1_7_out_E_noc3_yummy;
wire tile_1_7_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_2_7_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_2_7_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_2_7_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_2_7_out_W_noc1_data;
wire tile_2_7_out_N_noc1_valid;
wire tile_2_7_out_S_noc1_valid;
wire tile_2_7_out_E_noc1_valid;
wire tile_2_7_out_W_noc1_valid;
wire tile_2_7_out_N_noc1_yummy;
wire tile_2_7_out_S_noc1_yummy;
wire tile_2_7_out_E_noc1_yummy;
wire tile_2_7_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_2_7_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_2_7_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_2_7_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_2_7_out_W_noc2_data;
wire tile_2_7_out_N_noc2_valid;
wire tile_2_7_out_S_noc2_valid;
wire tile_2_7_out_E_noc2_valid;
wire tile_2_7_out_W_noc2_valid;
wire tile_2_7_out_N_noc2_yummy;
wire tile_2_7_out_S_noc2_yummy;
wire tile_2_7_out_E_noc2_yummy;
wire tile_2_7_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_2_7_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_2_7_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_2_7_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_2_7_out_W_noc3_data;
wire tile_2_7_out_N_noc3_valid;
wire tile_2_7_out_S_noc3_valid;
wire tile_2_7_out_E_noc3_valid;
wire tile_2_7_out_W_noc3_valid;
wire tile_2_7_out_N_noc3_yummy;
wire tile_2_7_out_S_noc3_yummy;
wire tile_2_7_out_E_noc3_yummy;
wire tile_2_7_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_3_7_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_3_7_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_3_7_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_3_7_out_W_noc1_data;
wire tile_3_7_out_N_noc1_valid;
wire tile_3_7_out_S_noc1_valid;
wire tile_3_7_out_E_noc1_valid;
wire tile_3_7_out_W_noc1_valid;
wire tile_3_7_out_N_noc1_yummy;
wire tile_3_7_out_S_noc1_yummy;
wire tile_3_7_out_E_noc1_yummy;
wire tile_3_7_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_3_7_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_3_7_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_3_7_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_3_7_out_W_noc2_data;
wire tile_3_7_out_N_noc2_valid;
wire tile_3_7_out_S_noc2_valid;
wire tile_3_7_out_E_noc2_valid;
wire tile_3_7_out_W_noc2_valid;
wire tile_3_7_out_N_noc2_yummy;
wire tile_3_7_out_S_noc2_yummy;
wire tile_3_7_out_E_noc2_yummy;
wire tile_3_7_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_3_7_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_3_7_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_3_7_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_3_7_out_W_noc3_data;
wire tile_3_7_out_N_noc3_valid;
wire tile_3_7_out_S_noc3_valid;
wire tile_3_7_out_E_noc3_valid;
wire tile_3_7_out_W_noc3_valid;
wire tile_3_7_out_N_noc3_yummy;
wire tile_3_7_out_S_noc3_yummy;
wire tile_3_7_out_E_noc3_yummy;
wire tile_3_7_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_4_7_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_4_7_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_4_7_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_4_7_out_W_noc1_data;
wire tile_4_7_out_N_noc1_valid;
wire tile_4_7_out_S_noc1_valid;
wire tile_4_7_out_E_noc1_valid;
wire tile_4_7_out_W_noc1_valid;
wire tile_4_7_out_N_noc1_yummy;
wire tile_4_7_out_S_noc1_yummy;
wire tile_4_7_out_E_noc1_yummy;
wire tile_4_7_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_4_7_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_4_7_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_4_7_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_4_7_out_W_noc2_data;
wire tile_4_7_out_N_noc2_valid;
wire tile_4_7_out_S_noc2_valid;
wire tile_4_7_out_E_noc2_valid;
wire tile_4_7_out_W_noc2_valid;
wire tile_4_7_out_N_noc2_yummy;
wire tile_4_7_out_S_noc2_yummy;
wire tile_4_7_out_E_noc2_yummy;
wire tile_4_7_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_4_7_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_4_7_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_4_7_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_4_7_out_W_noc3_data;
wire tile_4_7_out_N_noc3_valid;
wire tile_4_7_out_S_noc3_valid;
wire tile_4_7_out_E_noc3_valid;
wire tile_4_7_out_W_noc3_valid;
wire tile_4_7_out_N_noc3_yummy;
wire tile_4_7_out_S_noc3_yummy;
wire tile_4_7_out_E_noc3_yummy;
wire tile_4_7_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_5_7_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_5_7_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_5_7_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_5_7_out_W_noc1_data;
wire tile_5_7_out_N_noc1_valid;
wire tile_5_7_out_S_noc1_valid;
wire tile_5_7_out_E_noc1_valid;
wire tile_5_7_out_W_noc1_valid;
wire tile_5_7_out_N_noc1_yummy;
wire tile_5_7_out_S_noc1_yummy;
wire tile_5_7_out_E_noc1_yummy;
wire tile_5_7_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_5_7_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_5_7_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_5_7_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_5_7_out_W_noc2_data;
wire tile_5_7_out_N_noc2_valid;
wire tile_5_7_out_S_noc2_valid;
wire tile_5_7_out_E_noc2_valid;
wire tile_5_7_out_W_noc2_valid;
wire tile_5_7_out_N_noc2_yummy;
wire tile_5_7_out_S_noc2_yummy;
wire tile_5_7_out_E_noc2_yummy;
wire tile_5_7_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_5_7_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_5_7_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_5_7_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_5_7_out_W_noc3_data;
wire tile_5_7_out_N_noc3_valid;
wire tile_5_7_out_S_noc3_valid;
wire tile_5_7_out_E_noc3_valid;
wire tile_5_7_out_W_noc3_valid;
wire tile_5_7_out_N_noc3_yummy;
wire tile_5_7_out_S_noc3_yummy;
wire tile_5_7_out_E_noc3_yummy;
wire tile_5_7_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_6_7_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_6_7_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_6_7_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_6_7_out_W_noc1_data;
wire tile_6_7_out_N_noc1_valid;
wire tile_6_7_out_S_noc1_valid;
wire tile_6_7_out_E_noc1_valid;
wire tile_6_7_out_W_noc1_valid;
wire tile_6_7_out_N_noc1_yummy;
wire tile_6_7_out_S_noc1_yummy;
wire tile_6_7_out_E_noc1_yummy;
wire tile_6_7_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_6_7_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_6_7_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_6_7_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_6_7_out_W_noc2_data;
wire tile_6_7_out_N_noc2_valid;
wire tile_6_7_out_S_noc2_valid;
wire tile_6_7_out_E_noc2_valid;
wire tile_6_7_out_W_noc2_valid;
wire tile_6_7_out_N_noc2_yummy;
wire tile_6_7_out_S_noc2_yummy;
wire tile_6_7_out_E_noc2_yummy;
wire tile_6_7_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_6_7_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_6_7_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_6_7_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_6_7_out_W_noc3_data;
wire tile_6_7_out_N_noc3_valid;
wire tile_6_7_out_S_noc3_valid;
wire tile_6_7_out_E_noc3_valid;
wire tile_6_7_out_W_noc3_valid;
wire tile_6_7_out_N_noc3_yummy;
wire tile_6_7_out_S_noc3_yummy;
wire tile_6_7_out_E_noc3_yummy;
wire tile_6_7_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_7_7_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_7_7_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_7_7_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_7_7_out_W_noc1_data;
wire tile_7_7_out_N_noc1_valid;
wire tile_7_7_out_S_noc1_valid;
wire tile_7_7_out_E_noc1_valid;
wire tile_7_7_out_W_noc1_valid;
wire tile_7_7_out_N_noc1_yummy;
wire tile_7_7_out_S_noc1_yummy;
wire tile_7_7_out_E_noc1_yummy;
wire tile_7_7_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_7_7_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_7_7_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_7_7_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_7_7_out_W_noc2_data;
wire tile_7_7_out_N_noc2_valid;
wire tile_7_7_out_S_noc2_valid;
wire tile_7_7_out_E_noc2_valid;
wire tile_7_7_out_W_noc2_valid;
wire tile_7_7_out_N_noc2_yummy;
wire tile_7_7_out_S_noc2_yummy;
wire tile_7_7_out_E_noc2_yummy;
wire tile_7_7_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_7_7_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_7_7_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_7_7_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_7_7_out_W_noc3_data;
wire tile_7_7_out_N_noc3_valid;
wire tile_7_7_out_S_noc3_valid;
wire tile_7_7_out_E_noc3_valid;
wire tile_7_7_out_W_noc3_valid;
wire tile_7_7_out_N_noc3_yummy;
wire tile_7_7_out_S_noc3_yummy;
wire tile_7_7_out_E_noc3_yummy;
wire tile_7_7_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_8_7_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_8_7_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_8_7_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_8_7_out_W_noc1_data;
wire tile_8_7_out_N_noc1_valid;
wire tile_8_7_out_S_noc1_valid;
wire tile_8_7_out_E_noc1_valid;
wire tile_8_7_out_W_noc1_valid;
wire tile_8_7_out_N_noc1_yummy;
wire tile_8_7_out_S_noc1_yummy;
wire tile_8_7_out_E_noc1_yummy;
wire tile_8_7_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_8_7_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_8_7_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_8_7_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_8_7_out_W_noc2_data;
wire tile_8_7_out_N_noc2_valid;
wire tile_8_7_out_S_noc2_valid;
wire tile_8_7_out_E_noc2_valid;
wire tile_8_7_out_W_noc2_valid;
wire tile_8_7_out_N_noc2_yummy;
wire tile_8_7_out_S_noc2_yummy;
wire tile_8_7_out_E_noc2_yummy;
wire tile_8_7_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_8_7_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_8_7_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_8_7_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_8_7_out_W_noc3_data;
wire tile_8_7_out_N_noc3_valid;
wire tile_8_7_out_S_noc3_valid;
wire tile_8_7_out_E_noc3_valid;
wire tile_8_7_out_W_noc3_valid;
wire tile_8_7_out_N_noc3_yummy;
wire tile_8_7_out_S_noc3_yummy;
wire tile_8_7_out_E_noc3_yummy;
wire tile_8_7_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_9_7_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_9_7_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_9_7_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_9_7_out_W_noc1_data;
wire tile_9_7_out_N_noc1_valid;
wire tile_9_7_out_S_noc1_valid;
wire tile_9_7_out_E_noc1_valid;
wire tile_9_7_out_W_noc1_valid;
wire tile_9_7_out_N_noc1_yummy;
wire tile_9_7_out_S_noc1_yummy;
wire tile_9_7_out_E_noc1_yummy;
wire tile_9_7_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_9_7_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_9_7_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_9_7_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_9_7_out_W_noc2_data;
wire tile_9_7_out_N_noc2_valid;
wire tile_9_7_out_S_noc2_valid;
wire tile_9_7_out_E_noc2_valid;
wire tile_9_7_out_W_noc2_valid;
wire tile_9_7_out_N_noc2_yummy;
wire tile_9_7_out_S_noc2_yummy;
wire tile_9_7_out_E_noc2_yummy;
wire tile_9_7_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_9_7_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_9_7_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_9_7_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_9_7_out_W_noc3_data;
wire tile_9_7_out_N_noc3_valid;
wire tile_9_7_out_S_noc3_valid;
wire tile_9_7_out_E_noc3_valid;
wire tile_9_7_out_W_noc3_valid;
wire tile_9_7_out_N_noc3_yummy;
wire tile_9_7_out_S_noc3_yummy;
wire tile_9_7_out_E_noc3_yummy;
wire tile_9_7_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_10_7_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_10_7_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_10_7_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_10_7_out_W_noc1_data;
wire tile_10_7_out_N_noc1_valid;
wire tile_10_7_out_S_noc1_valid;
wire tile_10_7_out_E_noc1_valid;
wire tile_10_7_out_W_noc1_valid;
wire tile_10_7_out_N_noc1_yummy;
wire tile_10_7_out_S_noc1_yummy;
wire tile_10_7_out_E_noc1_yummy;
wire tile_10_7_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_10_7_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_10_7_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_10_7_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_10_7_out_W_noc2_data;
wire tile_10_7_out_N_noc2_valid;
wire tile_10_7_out_S_noc2_valid;
wire tile_10_7_out_E_noc2_valid;
wire tile_10_7_out_W_noc2_valid;
wire tile_10_7_out_N_noc2_yummy;
wire tile_10_7_out_S_noc2_yummy;
wire tile_10_7_out_E_noc2_yummy;
wire tile_10_7_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_10_7_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_10_7_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_10_7_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_10_7_out_W_noc3_data;
wire tile_10_7_out_N_noc3_valid;
wire tile_10_7_out_S_noc3_valid;
wire tile_10_7_out_E_noc3_valid;
wire tile_10_7_out_W_noc3_valid;
wire tile_10_7_out_N_noc3_yummy;
wire tile_10_7_out_S_noc3_yummy;
wire tile_10_7_out_E_noc3_yummy;
wire tile_10_7_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_11_7_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_11_7_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_11_7_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_11_7_out_W_noc1_data;
wire tile_11_7_out_N_noc1_valid;
wire tile_11_7_out_S_noc1_valid;
wire tile_11_7_out_E_noc1_valid;
wire tile_11_7_out_W_noc1_valid;
wire tile_11_7_out_N_noc1_yummy;
wire tile_11_7_out_S_noc1_yummy;
wire tile_11_7_out_E_noc1_yummy;
wire tile_11_7_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_11_7_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_11_7_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_11_7_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_11_7_out_W_noc2_data;
wire tile_11_7_out_N_noc2_valid;
wire tile_11_7_out_S_noc2_valid;
wire tile_11_7_out_E_noc2_valid;
wire tile_11_7_out_W_noc2_valid;
wire tile_11_7_out_N_noc2_yummy;
wire tile_11_7_out_S_noc2_yummy;
wire tile_11_7_out_E_noc2_yummy;
wire tile_11_7_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_11_7_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_11_7_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_11_7_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_11_7_out_W_noc3_data;
wire tile_11_7_out_N_noc3_valid;
wire tile_11_7_out_S_noc3_valid;
wire tile_11_7_out_E_noc3_valid;
wire tile_11_7_out_W_noc3_valid;
wire tile_11_7_out_N_noc3_yummy;
wire tile_11_7_out_S_noc3_yummy;
wire tile_11_7_out_E_noc3_yummy;
wire tile_11_7_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_12_7_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_12_7_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_12_7_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_12_7_out_W_noc1_data;
wire tile_12_7_out_N_noc1_valid;
wire tile_12_7_out_S_noc1_valid;
wire tile_12_7_out_E_noc1_valid;
wire tile_12_7_out_W_noc1_valid;
wire tile_12_7_out_N_noc1_yummy;
wire tile_12_7_out_S_noc1_yummy;
wire tile_12_7_out_E_noc1_yummy;
wire tile_12_7_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_12_7_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_12_7_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_12_7_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_12_7_out_W_noc2_data;
wire tile_12_7_out_N_noc2_valid;
wire tile_12_7_out_S_noc2_valid;
wire tile_12_7_out_E_noc2_valid;
wire tile_12_7_out_W_noc2_valid;
wire tile_12_7_out_N_noc2_yummy;
wire tile_12_7_out_S_noc2_yummy;
wire tile_12_7_out_E_noc2_yummy;
wire tile_12_7_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_12_7_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_12_7_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_12_7_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_12_7_out_W_noc3_data;
wire tile_12_7_out_N_noc3_valid;
wire tile_12_7_out_S_noc3_valid;
wire tile_12_7_out_E_noc3_valid;
wire tile_12_7_out_W_noc3_valid;
wire tile_12_7_out_N_noc3_yummy;
wire tile_12_7_out_S_noc3_yummy;
wire tile_12_7_out_E_noc3_yummy;
wire tile_12_7_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_13_7_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_13_7_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_13_7_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_13_7_out_W_noc1_data;
wire tile_13_7_out_N_noc1_valid;
wire tile_13_7_out_S_noc1_valid;
wire tile_13_7_out_E_noc1_valid;
wire tile_13_7_out_W_noc1_valid;
wire tile_13_7_out_N_noc1_yummy;
wire tile_13_7_out_S_noc1_yummy;
wire tile_13_7_out_E_noc1_yummy;
wire tile_13_7_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_13_7_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_13_7_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_13_7_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_13_7_out_W_noc2_data;
wire tile_13_7_out_N_noc2_valid;
wire tile_13_7_out_S_noc2_valid;
wire tile_13_7_out_E_noc2_valid;
wire tile_13_7_out_W_noc2_valid;
wire tile_13_7_out_N_noc2_yummy;
wire tile_13_7_out_S_noc2_yummy;
wire tile_13_7_out_E_noc2_yummy;
wire tile_13_7_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_13_7_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_13_7_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_13_7_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_13_7_out_W_noc3_data;
wire tile_13_7_out_N_noc3_valid;
wire tile_13_7_out_S_noc3_valid;
wire tile_13_7_out_E_noc3_valid;
wire tile_13_7_out_W_noc3_valid;
wire tile_13_7_out_N_noc3_yummy;
wire tile_13_7_out_S_noc3_yummy;
wire tile_13_7_out_E_noc3_yummy;
wire tile_13_7_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_14_7_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_14_7_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_14_7_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_14_7_out_W_noc1_data;
wire tile_14_7_out_N_noc1_valid;
wire tile_14_7_out_S_noc1_valid;
wire tile_14_7_out_E_noc1_valid;
wire tile_14_7_out_W_noc1_valid;
wire tile_14_7_out_N_noc1_yummy;
wire tile_14_7_out_S_noc1_yummy;
wire tile_14_7_out_E_noc1_yummy;
wire tile_14_7_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_14_7_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_14_7_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_14_7_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_14_7_out_W_noc2_data;
wire tile_14_7_out_N_noc2_valid;
wire tile_14_7_out_S_noc2_valid;
wire tile_14_7_out_E_noc2_valid;
wire tile_14_7_out_W_noc2_valid;
wire tile_14_7_out_N_noc2_yummy;
wire tile_14_7_out_S_noc2_yummy;
wire tile_14_7_out_E_noc2_yummy;
wire tile_14_7_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_14_7_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_14_7_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_14_7_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_14_7_out_W_noc3_data;
wire tile_14_7_out_N_noc3_valid;
wire tile_14_7_out_S_noc3_valid;
wire tile_14_7_out_E_noc3_valid;
wire tile_14_7_out_W_noc3_valid;
wire tile_14_7_out_N_noc3_yummy;
wire tile_14_7_out_S_noc3_yummy;
wire tile_14_7_out_E_noc3_yummy;
wire tile_14_7_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_15_7_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_15_7_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_15_7_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_15_7_out_W_noc1_data;
wire tile_15_7_out_N_noc1_valid;
wire tile_15_7_out_S_noc1_valid;
wire tile_15_7_out_E_noc1_valid;
wire tile_15_7_out_W_noc1_valid;
wire tile_15_7_out_N_noc1_yummy;
wire tile_15_7_out_S_noc1_yummy;
wire tile_15_7_out_E_noc1_yummy;
wire tile_15_7_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_15_7_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_15_7_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_15_7_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_15_7_out_W_noc2_data;
wire tile_15_7_out_N_noc2_valid;
wire tile_15_7_out_S_noc2_valid;
wire tile_15_7_out_E_noc2_valid;
wire tile_15_7_out_W_noc2_valid;
wire tile_15_7_out_N_noc2_yummy;
wire tile_15_7_out_S_noc2_yummy;
wire tile_15_7_out_E_noc2_yummy;
wire tile_15_7_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_15_7_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_15_7_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_15_7_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_15_7_out_W_noc3_data;
wire tile_15_7_out_N_noc3_valid;
wire tile_15_7_out_S_noc3_valid;
wire tile_15_7_out_E_noc3_valid;
wire tile_15_7_out_W_noc3_valid;
wire tile_15_7_out_N_noc3_yummy;
wire tile_15_7_out_S_noc3_yummy;
wire tile_15_7_out_E_noc3_yummy;
wire tile_15_7_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_0_8_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_0_8_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_0_8_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_0_8_out_W_noc1_data;
wire tile_0_8_out_N_noc1_valid;
wire tile_0_8_out_S_noc1_valid;
wire tile_0_8_out_E_noc1_valid;
wire tile_0_8_out_W_noc1_valid;
wire tile_0_8_out_N_noc1_yummy;
wire tile_0_8_out_S_noc1_yummy;
wire tile_0_8_out_E_noc1_yummy;
wire tile_0_8_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_0_8_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_0_8_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_0_8_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_0_8_out_W_noc2_data;
wire tile_0_8_out_N_noc2_valid;
wire tile_0_8_out_S_noc2_valid;
wire tile_0_8_out_E_noc2_valid;
wire tile_0_8_out_W_noc2_valid;
wire tile_0_8_out_N_noc2_yummy;
wire tile_0_8_out_S_noc2_yummy;
wire tile_0_8_out_E_noc2_yummy;
wire tile_0_8_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_0_8_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_0_8_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_0_8_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_0_8_out_W_noc3_data;
wire tile_0_8_out_N_noc3_valid;
wire tile_0_8_out_S_noc3_valid;
wire tile_0_8_out_E_noc3_valid;
wire tile_0_8_out_W_noc3_valid;
wire tile_0_8_out_N_noc3_yummy;
wire tile_0_8_out_S_noc3_yummy;
wire tile_0_8_out_E_noc3_yummy;
wire tile_0_8_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_1_8_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_1_8_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_1_8_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_1_8_out_W_noc1_data;
wire tile_1_8_out_N_noc1_valid;
wire tile_1_8_out_S_noc1_valid;
wire tile_1_8_out_E_noc1_valid;
wire tile_1_8_out_W_noc1_valid;
wire tile_1_8_out_N_noc1_yummy;
wire tile_1_8_out_S_noc1_yummy;
wire tile_1_8_out_E_noc1_yummy;
wire tile_1_8_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_1_8_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_1_8_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_1_8_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_1_8_out_W_noc2_data;
wire tile_1_8_out_N_noc2_valid;
wire tile_1_8_out_S_noc2_valid;
wire tile_1_8_out_E_noc2_valid;
wire tile_1_8_out_W_noc2_valid;
wire tile_1_8_out_N_noc2_yummy;
wire tile_1_8_out_S_noc2_yummy;
wire tile_1_8_out_E_noc2_yummy;
wire tile_1_8_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_1_8_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_1_8_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_1_8_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_1_8_out_W_noc3_data;
wire tile_1_8_out_N_noc3_valid;
wire tile_1_8_out_S_noc3_valid;
wire tile_1_8_out_E_noc3_valid;
wire tile_1_8_out_W_noc3_valid;
wire tile_1_8_out_N_noc3_yummy;
wire tile_1_8_out_S_noc3_yummy;
wire tile_1_8_out_E_noc3_yummy;
wire tile_1_8_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_2_8_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_2_8_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_2_8_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_2_8_out_W_noc1_data;
wire tile_2_8_out_N_noc1_valid;
wire tile_2_8_out_S_noc1_valid;
wire tile_2_8_out_E_noc1_valid;
wire tile_2_8_out_W_noc1_valid;
wire tile_2_8_out_N_noc1_yummy;
wire tile_2_8_out_S_noc1_yummy;
wire tile_2_8_out_E_noc1_yummy;
wire tile_2_8_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_2_8_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_2_8_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_2_8_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_2_8_out_W_noc2_data;
wire tile_2_8_out_N_noc2_valid;
wire tile_2_8_out_S_noc2_valid;
wire tile_2_8_out_E_noc2_valid;
wire tile_2_8_out_W_noc2_valid;
wire tile_2_8_out_N_noc2_yummy;
wire tile_2_8_out_S_noc2_yummy;
wire tile_2_8_out_E_noc2_yummy;
wire tile_2_8_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_2_8_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_2_8_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_2_8_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_2_8_out_W_noc3_data;
wire tile_2_8_out_N_noc3_valid;
wire tile_2_8_out_S_noc3_valid;
wire tile_2_8_out_E_noc3_valid;
wire tile_2_8_out_W_noc3_valid;
wire tile_2_8_out_N_noc3_yummy;
wire tile_2_8_out_S_noc3_yummy;
wire tile_2_8_out_E_noc3_yummy;
wire tile_2_8_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_3_8_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_3_8_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_3_8_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_3_8_out_W_noc1_data;
wire tile_3_8_out_N_noc1_valid;
wire tile_3_8_out_S_noc1_valid;
wire tile_3_8_out_E_noc1_valid;
wire tile_3_8_out_W_noc1_valid;
wire tile_3_8_out_N_noc1_yummy;
wire tile_3_8_out_S_noc1_yummy;
wire tile_3_8_out_E_noc1_yummy;
wire tile_3_8_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_3_8_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_3_8_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_3_8_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_3_8_out_W_noc2_data;
wire tile_3_8_out_N_noc2_valid;
wire tile_3_8_out_S_noc2_valid;
wire tile_3_8_out_E_noc2_valid;
wire tile_3_8_out_W_noc2_valid;
wire tile_3_8_out_N_noc2_yummy;
wire tile_3_8_out_S_noc2_yummy;
wire tile_3_8_out_E_noc2_yummy;
wire tile_3_8_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_3_8_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_3_8_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_3_8_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_3_8_out_W_noc3_data;
wire tile_3_8_out_N_noc3_valid;
wire tile_3_8_out_S_noc3_valid;
wire tile_3_8_out_E_noc3_valid;
wire tile_3_8_out_W_noc3_valid;
wire tile_3_8_out_N_noc3_yummy;
wire tile_3_8_out_S_noc3_yummy;
wire tile_3_8_out_E_noc3_yummy;
wire tile_3_8_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_4_8_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_4_8_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_4_8_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_4_8_out_W_noc1_data;
wire tile_4_8_out_N_noc1_valid;
wire tile_4_8_out_S_noc1_valid;
wire tile_4_8_out_E_noc1_valid;
wire tile_4_8_out_W_noc1_valid;
wire tile_4_8_out_N_noc1_yummy;
wire tile_4_8_out_S_noc1_yummy;
wire tile_4_8_out_E_noc1_yummy;
wire tile_4_8_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_4_8_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_4_8_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_4_8_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_4_8_out_W_noc2_data;
wire tile_4_8_out_N_noc2_valid;
wire tile_4_8_out_S_noc2_valid;
wire tile_4_8_out_E_noc2_valid;
wire tile_4_8_out_W_noc2_valid;
wire tile_4_8_out_N_noc2_yummy;
wire tile_4_8_out_S_noc2_yummy;
wire tile_4_8_out_E_noc2_yummy;
wire tile_4_8_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_4_8_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_4_8_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_4_8_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_4_8_out_W_noc3_data;
wire tile_4_8_out_N_noc3_valid;
wire tile_4_8_out_S_noc3_valid;
wire tile_4_8_out_E_noc3_valid;
wire tile_4_8_out_W_noc3_valid;
wire tile_4_8_out_N_noc3_yummy;
wire tile_4_8_out_S_noc3_yummy;
wire tile_4_8_out_E_noc3_yummy;
wire tile_4_8_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_5_8_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_5_8_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_5_8_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_5_8_out_W_noc1_data;
wire tile_5_8_out_N_noc1_valid;
wire tile_5_8_out_S_noc1_valid;
wire tile_5_8_out_E_noc1_valid;
wire tile_5_8_out_W_noc1_valid;
wire tile_5_8_out_N_noc1_yummy;
wire tile_5_8_out_S_noc1_yummy;
wire tile_5_8_out_E_noc1_yummy;
wire tile_5_8_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_5_8_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_5_8_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_5_8_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_5_8_out_W_noc2_data;
wire tile_5_8_out_N_noc2_valid;
wire tile_5_8_out_S_noc2_valid;
wire tile_5_8_out_E_noc2_valid;
wire tile_5_8_out_W_noc2_valid;
wire tile_5_8_out_N_noc2_yummy;
wire tile_5_8_out_S_noc2_yummy;
wire tile_5_8_out_E_noc2_yummy;
wire tile_5_8_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_5_8_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_5_8_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_5_8_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_5_8_out_W_noc3_data;
wire tile_5_8_out_N_noc3_valid;
wire tile_5_8_out_S_noc3_valid;
wire tile_5_8_out_E_noc3_valid;
wire tile_5_8_out_W_noc3_valid;
wire tile_5_8_out_N_noc3_yummy;
wire tile_5_8_out_S_noc3_yummy;
wire tile_5_8_out_E_noc3_yummy;
wire tile_5_8_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_6_8_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_6_8_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_6_8_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_6_8_out_W_noc1_data;
wire tile_6_8_out_N_noc1_valid;
wire tile_6_8_out_S_noc1_valid;
wire tile_6_8_out_E_noc1_valid;
wire tile_6_8_out_W_noc1_valid;
wire tile_6_8_out_N_noc1_yummy;
wire tile_6_8_out_S_noc1_yummy;
wire tile_6_8_out_E_noc1_yummy;
wire tile_6_8_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_6_8_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_6_8_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_6_8_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_6_8_out_W_noc2_data;
wire tile_6_8_out_N_noc2_valid;
wire tile_6_8_out_S_noc2_valid;
wire tile_6_8_out_E_noc2_valid;
wire tile_6_8_out_W_noc2_valid;
wire tile_6_8_out_N_noc2_yummy;
wire tile_6_8_out_S_noc2_yummy;
wire tile_6_8_out_E_noc2_yummy;
wire tile_6_8_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_6_8_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_6_8_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_6_8_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_6_8_out_W_noc3_data;
wire tile_6_8_out_N_noc3_valid;
wire tile_6_8_out_S_noc3_valid;
wire tile_6_8_out_E_noc3_valid;
wire tile_6_8_out_W_noc3_valid;
wire tile_6_8_out_N_noc3_yummy;
wire tile_6_8_out_S_noc3_yummy;
wire tile_6_8_out_E_noc3_yummy;
wire tile_6_8_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_7_8_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_7_8_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_7_8_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_7_8_out_W_noc1_data;
wire tile_7_8_out_N_noc1_valid;
wire tile_7_8_out_S_noc1_valid;
wire tile_7_8_out_E_noc1_valid;
wire tile_7_8_out_W_noc1_valid;
wire tile_7_8_out_N_noc1_yummy;
wire tile_7_8_out_S_noc1_yummy;
wire tile_7_8_out_E_noc1_yummy;
wire tile_7_8_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_7_8_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_7_8_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_7_8_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_7_8_out_W_noc2_data;
wire tile_7_8_out_N_noc2_valid;
wire tile_7_8_out_S_noc2_valid;
wire tile_7_8_out_E_noc2_valid;
wire tile_7_8_out_W_noc2_valid;
wire tile_7_8_out_N_noc2_yummy;
wire tile_7_8_out_S_noc2_yummy;
wire tile_7_8_out_E_noc2_yummy;
wire tile_7_8_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_7_8_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_7_8_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_7_8_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_7_8_out_W_noc3_data;
wire tile_7_8_out_N_noc3_valid;
wire tile_7_8_out_S_noc3_valid;
wire tile_7_8_out_E_noc3_valid;
wire tile_7_8_out_W_noc3_valid;
wire tile_7_8_out_N_noc3_yummy;
wire tile_7_8_out_S_noc3_yummy;
wire tile_7_8_out_E_noc3_yummy;
wire tile_7_8_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_8_8_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_8_8_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_8_8_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_8_8_out_W_noc1_data;
wire tile_8_8_out_N_noc1_valid;
wire tile_8_8_out_S_noc1_valid;
wire tile_8_8_out_E_noc1_valid;
wire tile_8_8_out_W_noc1_valid;
wire tile_8_8_out_N_noc1_yummy;
wire tile_8_8_out_S_noc1_yummy;
wire tile_8_8_out_E_noc1_yummy;
wire tile_8_8_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_8_8_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_8_8_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_8_8_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_8_8_out_W_noc2_data;
wire tile_8_8_out_N_noc2_valid;
wire tile_8_8_out_S_noc2_valid;
wire tile_8_8_out_E_noc2_valid;
wire tile_8_8_out_W_noc2_valid;
wire tile_8_8_out_N_noc2_yummy;
wire tile_8_8_out_S_noc2_yummy;
wire tile_8_8_out_E_noc2_yummy;
wire tile_8_8_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_8_8_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_8_8_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_8_8_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_8_8_out_W_noc3_data;
wire tile_8_8_out_N_noc3_valid;
wire tile_8_8_out_S_noc3_valid;
wire tile_8_8_out_E_noc3_valid;
wire tile_8_8_out_W_noc3_valid;
wire tile_8_8_out_N_noc3_yummy;
wire tile_8_8_out_S_noc3_yummy;
wire tile_8_8_out_E_noc3_yummy;
wire tile_8_8_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_9_8_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_9_8_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_9_8_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_9_8_out_W_noc1_data;
wire tile_9_8_out_N_noc1_valid;
wire tile_9_8_out_S_noc1_valid;
wire tile_9_8_out_E_noc1_valid;
wire tile_9_8_out_W_noc1_valid;
wire tile_9_8_out_N_noc1_yummy;
wire tile_9_8_out_S_noc1_yummy;
wire tile_9_8_out_E_noc1_yummy;
wire tile_9_8_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_9_8_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_9_8_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_9_8_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_9_8_out_W_noc2_data;
wire tile_9_8_out_N_noc2_valid;
wire tile_9_8_out_S_noc2_valid;
wire tile_9_8_out_E_noc2_valid;
wire tile_9_8_out_W_noc2_valid;
wire tile_9_8_out_N_noc2_yummy;
wire tile_9_8_out_S_noc2_yummy;
wire tile_9_8_out_E_noc2_yummy;
wire tile_9_8_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_9_8_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_9_8_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_9_8_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_9_8_out_W_noc3_data;
wire tile_9_8_out_N_noc3_valid;
wire tile_9_8_out_S_noc3_valid;
wire tile_9_8_out_E_noc3_valid;
wire tile_9_8_out_W_noc3_valid;
wire tile_9_8_out_N_noc3_yummy;
wire tile_9_8_out_S_noc3_yummy;
wire tile_9_8_out_E_noc3_yummy;
wire tile_9_8_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_10_8_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_10_8_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_10_8_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_10_8_out_W_noc1_data;
wire tile_10_8_out_N_noc1_valid;
wire tile_10_8_out_S_noc1_valid;
wire tile_10_8_out_E_noc1_valid;
wire tile_10_8_out_W_noc1_valid;
wire tile_10_8_out_N_noc1_yummy;
wire tile_10_8_out_S_noc1_yummy;
wire tile_10_8_out_E_noc1_yummy;
wire tile_10_8_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_10_8_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_10_8_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_10_8_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_10_8_out_W_noc2_data;
wire tile_10_8_out_N_noc2_valid;
wire tile_10_8_out_S_noc2_valid;
wire tile_10_8_out_E_noc2_valid;
wire tile_10_8_out_W_noc2_valid;
wire tile_10_8_out_N_noc2_yummy;
wire tile_10_8_out_S_noc2_yummy;
wire tile_10_8_out_E_noc2_yummy;
wire tile_10_8_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_10_8_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_10_8_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_10_8_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_10_8_out_W_noc3_data;
wire tile_10_8_out_N_noc3_valid;
wire tile_10_8_out_S_noc3_valid;
wire tile_10_8_out_E_noc3_valid;
wire tile_10_8_out_W_noc3_valid;
wire tile_10_8_out_N_noc3_yummy;
wire tile_10_8_out_S_noc3_yummy;
wire tile_10_8_out_E_noc3_yummy;
wire tile_10_8_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_11_8_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_11_8_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_11_8_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_11_8_out_W_noc1_data;
wire tile_11_8_out_N_noc1_valid;
wire tile_11_8_out_S_noc1_valid;
wire tile_11_8_out_E_noc1_valid;
wire tile_11_8_out_W_noc1_valid;
wire tile_11_8_out_N_noc1_yummy;
wire tile_11_8_out_S_noc1_yummy;
wire tile_11_8_out_E_noc1_yummy;
wire tile_11_8_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_11_8_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_11_8_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_11_8_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_11_8_out_W_noc2_data;
wire tile_11_8_out_N_noc2_valid;
wire tile_11_8_out_S_noc2_valid;
wire tile_11_8_out_E_noc2_valid;
wire tile_11_8_out_W_noc2_valid;
wire tile_11_8_out_N_noc2_yummy;
wire tile_11_8_out_S_noc2_yummy;
wire tile_11_8_out_E_noc2_yummy;
wire tile_11_8_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_11_8_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_11_8_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_11_8_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_11_8_out_W_noc3_data;
wire tile_11_8_out_N_noc3_valid;
wire tile_11_8_out_S_noc3_valid;
wire tile_11_8_out_E_noc3_valid;
wire tile_11_8_out_W_noc3_valid;
wire tile_11_8_out_N_noc3_yummy;
wire tile_11_8_out_S_noc3_yummy;
wire tile_11_8_out_E_noc3_yummy;
wire tile_11_8_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_12_8_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_12_8_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_12_8_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_12_8_out_W_noc1_data;
wire tile_12_8_out_N_noc1_valid;
wire tile_12_8_out_S_noc1_valid;
wire tile_12_8_out_E_noc1_valid;
wire tile_12_8_out_W_noc1_valid;
wire tile_12_8_out_N_noc1_yummy;
wire tile_12_8_out_S_noc1_yummy;
wire tile_12_8_out_E_noc1_yummy;
wire tile_12_8_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_12_8_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_12_8_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_12_8_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_12_8_out_W_noc2_data;
wire tile_12_8_out_N_noc2_valid;
wire tile_12_8_out_S_noc2_valid;
wire tile_12_8_out_E_noc2_valid;
wire tile_12_8_out_W_noc2_valid;
wire tile_12_8_out_N_noc2_yummy;
wire tile_12_8_out_S_noc2_yummy;
wire tile_12_8_out_E_noc2_yummy;
wire tile_12_8_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_12_8_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_12_8_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_12_8_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_12_8_out_W_noc3_data;
wire tile_12_8_out_N_noc3_valid;
wire tile_12_8_out_S_noc3_valid;
wire tile_12_8_out_E_noc3_valid;
wire tile_12_8_out_W_noc3_valid;
wire tile_12_8_out_N_noc3_yummy;
wire tile_12_8_out_S_noc3_yummy;
wire tile_12_8_out_E_noc3_yummy;
wire tile_12_8_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_13_8_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_13_8_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_13_8_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_13_8_out_W_noc1_data;
wire tile_13_8_out_N_noc1_valid;
wire tile_13_8_out_S_noc1_valid;
wire tile_13_8_out_E_noc1_valid;
wire tile_13_8_out_W_noc1_valid;
wire tile_13_8_out_N_noc1_yummy;
wire tile_13_8_out_S_noc1_yummy;
wire tile_13_8_out_E_noc1_yummy;
wire tile_13_8_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_13_8_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_13_8_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_13_8_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_13_8_out_W_noc2_data;
wire tile_13_8_out_N_noc2_valid;
wire tile_13_8_out_S_noc2_valid;
wire tile_13_8_out_E_noc2_valid;
wire tile_13_8_out_W_noc2_valid;
wire tile_13_8_out_N_noc2_yummy;
wire tile_13_8_out_S_noc2_yummy;
wire tile_13_8_out_E_noc2_yummy;
wire tile_13_8_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_13_8_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_13_8_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_13_8_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_13_8_out_W_noc3_data;
wire tile_13_8_out_N_noc3_valid;
wire tile_13_8_out_S_noc3_valid;
wire tile_13_8_out_E_noc3_valid;
wire tile_13_8_out_W_noc3_valid;
wire tile_13_8_out_N_noc3_yummy;
wire tile_13_8_out_S_noc3_yummy;
wire tile_13_8_out_E_noc3_yummy;
wire tile_13_8_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_14_8_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_14_8_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_14_8_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_14_8_out_W_noc1_data;
wire tile_14_8_out_N_noc1_valid;
wire tile_14_8_out_S_noc1_valid;
wire tile_14_8_out_E_noc1_valid;
wire tile_14_8_out_W_noc1_valid;
wire tile_14_8_out_N_noc1_yummy;
wire tile_14_8_out_S_noc1_yummy;
wire tile_14_8_out_E_noc1_yummy;
wire tile_14_8_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_14_8_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_14_8_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_14_8_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_14_8_out_W_noc2_data;
wire tile_14_8_out_N_noc2_valid;
wire tile_14_8_out_S_noc2_valid;
wire tile_14_8_out_E_noc2_valid;
wire tile_14_8_out_W_noc2_valid;
wire tile_14_8_out_N_noc2_yummy;
wire tile_14_8_out_S_noc2_yummy;
wire tile_14_8_out_E_noc2_yummy;
wire tile_14_8_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_14_8_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_14_8_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_14_8_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_14_8_out_W_noc3_data;
wire tile_14_8_out_N_noc3_valid;
wire tile_14_8_out_S_noc3_valid;
wire tile_14_8_out_E_noc3_valid;
wire tile_14_8_out_W_noc3_valid;
wire tile_14_8_out_N_noc3_yummy;
wire tile_14_8_out_S_noc3_yummy;
wire tile_14_8_out_E_noc3_yummy;
wire tile_14_8_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_15_8_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_15_8_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_15_8_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_15_8_out_W_noc1_data;
wire tile_15_8_out_N_noc1_valid;
wire tile_15_8_out_S_noc1_valid;
wire tile_15_8_out_E_noc1_valid;
wire tile_15_8_out_W_noc1_valid;
wire tile_15_8_out_N_noc1_yummy;
wire tile_15_8_out_S_noc1_yummy;
wire tile_15_8_out_E_noc1_yummy;
wire tile_15_8_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_15_8_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_15_8_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_15_8_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_15_8_out_W_noc2_data;
wire tile_15_8_out_N_noc2_valid;
wire tile_15_8_out_S_noc2_valid;
wire tile_15_8_out_E_noc2_valid;
wire tile_15_8_out_W_noc2_valid;
wire tile_15_8_out_N_noc2_yummy;
wire tile_15_8_out_S_noc2_yummy;
wire tile_15_8_out_E_noc2_yummy;
wire tile_15_8_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_15_8_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_15_8_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_15_8_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_15_8_out_W_noc3_data;
wire tile_15_8_out_N_noc3_valid;
wire tile_15_8_out_S_noc3_valid;
wire tile_15_8_out_E_noc3_valid;
wire tile_15_8_out_W_noc3_valid;
wire tile_15_8_out_N_noc3_yummy;
wire tile_15_8_out_S_noc3_yummy;
wire tile_15_8_out_E_noc3_yummy;
wire tile_15_8_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_0_9_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_0_9_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_0_9_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_0_9_out_W_noc1_data;
wire tile_0_9_out_N_noc1_valid;
wire tile_0_9_out_S_noc1_valid;
wire tile_0_9_out_E_noc1_valid;
wire tile_0_9_out_W_noc1_valid;
wire tile_0_9_out_N_noc1_yummy;
wire tile_0_9_out_S_noc1_yummy;
wire tile_0_9_out_E_noc1_yummy;
wire tile_0_9_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_0_9_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_0_9_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_0_9_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_0_9_out_W_noc2_data;
wire tile_0_9_out_N_noc2_valid;
wire tile_0_9_out_S_noc2_valid;
wire tile_0_9_out_E_noc2_valid;
wire tile_0_9_out_W_noc2_valid;
wire tile_0_9_out_N_noc2_yummy;
wire tile_0_9_out_S_noc2_yummy;
wire tile_0_9_out_E_noc2_yummy;
wire tile_0_9_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_0_9_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_0_9_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_0_9_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_0_9_out_W_noc3_data;
wire tile_0_9_out_N_noc3_valid;
wire tile_0_9_out_S_noc3_valid;
wire tile_0_9_out_E_noc3_valid;
wire tile_0_9_out_W_noc3_valid;
wire tile_0_9_out_N_noc3_yummy;
wire tile_0_9_out_S_noc3_yummy;
wire tile_0_9_out_E_noc3_yummy;
wire tile_0_9_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_1_9_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_1_9_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_1_9_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_1_9_out_W_noc1_data;
wire tile_1_9_out_N_noc1_valid;
wire tile_1_9_out_S_noc1_valid;
wire tile_1_9_out_E_noc1_valid;
wire tile_1_9_out_W_noc1_valid;
wire tile_1_9_out_N_noc1_yummy;
wire tile_1_9_out_S_noc1_yummy;
wire tile_1_9_out_E_noc1_yummy;
wire tile_1_9_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_1_9_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_1_9_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_1_9_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_1_9_out_W_noc2_data;
wire tile_1_9_out_N_noc2_valid;
wire tile_1_9_out_S_noc2_valid;
wire tile_1_9_out_E_noc2_valid;
wire tile_1_9_out_W_noc2_valid;
wire tile_1_9_out_N_noc2_yummy;
wire tile_1_9_out_S_noc2_yummy;
wire tile_1_9_out_E_noc2_yummy;
wire tile_1_9_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_1_9_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_1_9_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_1_9_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_1_9_out_W_noc3_data;
wire tile_1_9_out_N_noc3_valid;
wire tile_1_9_out_S_noc3_valid;
wire tile_1_9_out_E_noc3_valid;
wire tile_1_9_out_W_noc3_valid;
wire tile_1_9_out_N_noc3_yummy;
wire tile_1_9_out_S_noc3_yummy;
wire tile_1_9_out_E_noc3_yummy;
wire tile_1_9_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_2_9_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_2_9_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_2_9_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_2_9_out_W_noc1_data;
wire tile_2_9_out_N_noc1_valid;
wire tile_2_9_out_S_noc1_valid;
wire tile_2_9_out_E_noc1_valid;
wire tile_2_9_out_W_noc1_valid;
wire tile_2_9_out_N_noc1_yummy;
wire tile_2_9_out_S_noc1_yummy;
wire tile_2_9_out_E_noc1_yummy;
wire tile_2_9_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_2_9_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_2_9_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_2_9_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_2_9_out_W_noc2_data;
wire tile_2_9_out_N_noc2_valid;
wire tile_2_9_out_S_noc2_valid;
wire tile_2_9_out_E_noc2_valid;
wire tile_2_9_out_W_noc2_valid;
wire tile_2_9_out_N_noc2_yummy;
wire tile_2_9_out_S_noc2_yummy;
wire tile_2_9_out_E_noc2_yummy;
wire tile_2_9_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_2_9_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_2_9_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_2_9_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_2_9_out_W_noc3_data;
wire tile_2_9_out_N_noc3_valid;
wire tile_2_9_out_S_noc3_valid;
wire tile_2_9_out_E_noc3_valid;
wire tile_2_9_out_W_noc3_valid;
wire tile_2_9_out_N_noc3_yummy;
wire tile_2_9_out_S_noc3_yummy;
wire tile_2_9_out_E_noc3_yummy;
wire tile_2_9_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_3_9_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_3_9_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_3_9_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_3_9_out_W_noc1_data;
wire tile_3_9_out_N_noc1_valid;
wire tile_3_9_out_S_noc1_valid;
wire tile_3_9_out_E_noc1_valid;
wire tile_3_9_out_W_noc1_valid;
wire tile_3_9_out_N_noc1_yummy;
wire tile_3_9_out_S_noc1_yummy;
wire tile_3_9_out_E_noc1_yummy;
wire tile_3_9_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_3_9_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_3_9_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_3_9_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_3_9_out_W_noc2_data;
wire tile_3_9_out_N_noc2_valid;
wire tile_3_9_out_S_noc2_valid;
wire tile_3_9_out_E_noc2_valid;
wire tile_3_9_out_W_noc2_valid;
wire tile_3_9_out_N_noc2_yummy;
wire tile_3_9_out_S_noc2_yummy;
wire tile_3_9_out_E_noc2_yummy;
wire tile_3_9_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_3_9_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_3_9_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_3_9_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_3_9_out_W_noc3_data;
wire tile_3_9_out_N_noc3_valid;
wire tile_3_9_out_S_noc3_valid;
wire tile_3_9_out_E_noc3_valid;
wire tile_3_9_out_W_noc3_valid;
wire tile_3_9_out_N_noc3_yummy;
wire tile_3_9_out_S_noc3_yummy;
wire tile_3_9_out_E_noc3_yummy;
wire tile_3_9_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_4_9_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_4_9_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_4_9_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_4_9_out_W_noc1_data;
wire tile_4_9_out_N_noc1_valid;
wire tile_4_9_out_S_noc1_valid;
wire tile_4_9_out_E_noc1_valid;
wire tile_4_9_out_W_noc1_valid;
wire tile_4_9_out_N_noc1_yummy;
wire tile_4_9_out_S_noc1_yummy;
wire tile_4_9_out_E_noc1_yummy;
wire tile_4_9_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_4_9_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_4_9_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_4_9_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_4_9_out_W_noc2_data;
wire tile_4_9_out_N_noc2_valid;
wire tile_4_9_out_S_noc2_valid;
wire tile_4_9_out_E_noc2_valid;
wire tile_4_9_out_W_noc2_valid;
wire tile_4_9_out_N_noc2_yummy;
wire tile_4_9_out_S_noc2_yummy;
wire tile_4_9_out_E_noc2_yummy;
wire tile_4_9_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_4_9_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_4_9_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_4_9_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_4_9_out_W_noc3_data;
wire tile_4_9_out_N_noc3_valid;
wire tile_4_9_out_S_noc3_valid;
wire tile_4_9_out_E_noc3_valid;
wire tile_4_9_out_W_noc3_valid;
wire tile_4_9_out_N_noc3_yummy;
wire tile_4_9_out_S_noc3_yummy;
wire tile_4_9_out_E_noc3_yummy;
wire tile_4_9_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_5_9_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_5_9_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_5_9_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_5_9_out_W_noc1_data;
wire tile_5_9_out_N_noc1_valid;
wire tile_5_9_out_S_noc1_valid;
wire tile_5_9_out_E_noc1_valid;
wire tile_5_9_out_W_noc1_valid;
wire tile_5_9_out_N_noc1_yummy;
wire tile_5_9_out_S_noc1_yummy;
wire tile_5_9_out_E_noc1_yummy;
wire tile_5_9_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_5_9_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_5_9_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_5_9_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_5_9_out_W_noc2_data;
wire tile_5_9_out_N_noc2_valid;
wire tile_5_9_out_S_noc2_valid;
wire tile_5_9_out_E_noc2_valid;
wire tile_5_9_out_W_noc2_valid;
wire tile_5_9_out_N_noc2_yummy;
wire tile_5_9_out_S_noc2_yummy;
wire tile_5_9_out_E_noc2_yummy;
wire tile_5_9_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_5_9_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_5_9_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_5_9_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_5_9_out_W_noc3_data;
wire tile_5_9_out_N_noc3_valid;
wire tile_5_9_out_S_noc3_valid;
wire tile_5_9_out_E_noc3_valid;
wire tile_5_9_out_W_noc3_valid;
wire tile_5_9_out_N_noc3_yummy;
wire tile_5_9_out_S_noc3_yummy;
wire tile_5_9_out_E_noc3_yummy;
wire tile_5_9_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_6_9_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_6_9_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_6_9_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_6_9_out_W_noc1_data;
wire tile_6_9_out_N_noc1_valid;
wire tile_6_9_out_S_noc1_valid;
wire tile_6_9_out_E_noc1_valid;
wire tile_6_9_out_W_noc1_valid;
wire tile_6_9_out_N_noc1_yummy;
wire tile_6_9_out_S_noc1_yummy;
wire tile_6_9_out_E_noc1_yummy;
wire tile_6_9_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_6_9_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_6_9_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_6_9_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_6_9_out_W_noc2_data;
wire tile_6_9_out_N_noc2_valid;
wire tile_6_9_out_S_noc2_valid;
wire tile_6_9_out_E_noc2_valid;
wire tile_6_9_out_W_noc2_valid;
wire tile_6_9_out_N_noc2_yummy;
wire tile_6_9_out_S_noc2_yummy;
wire tile_6_9_out_E_noc2_yummy;
wire tile_6_9_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_6_9_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_6_9_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_6_9_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_6_9_out_W_noc3_data;
wire tile_6_9_out_N_noc3_valid;
wire tile_6_9_out_S_noc3_valid;
wire tile_6_9_out_E_noc3_valid;
wire tile_6_9_out_W_noc3_valid;
wire tile_6_9_out_N_noc3_yummy;
wire tile_6_9_out_S_noc3_yummy;
wire tile_6_9_out_E_noc3_yummy;
wire tile_6_9_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_7_9_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_7_9_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_7_9_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_7_9_out_W_noc1_data;
wire tile_7_9_out_N_noc1_valid;
wire tile_7_9_out_S_noc1_valid;
wire tile_7_9_out_E_noc1_valid;
wire tile_7_9_out_W_noc1_valid;
wire tile_7_9_out_N_noc1_yummy;
wire tile_7_9_out_S_noc1_yummy;
wire tile_7_9_out_E_noc1_yummy;
wire tile_7_9_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_7_9_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_7_9_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_7_9_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_7_9_out_W_noc2_data;
wire tile_7_9_out_N_noc2_valid;
wire tile_7_9_out_S_noc2_valid;
wire tile_7_9_out_E_noc2_valid;
wire tile_7_9_out_W_noc2_valid;
wire tile_7_9_out_N_noc2_yummy;
wire tile_7_9_out_S_noc2_yummy;
wire tile_7_9_out_E_noc2_yummy;
wire tile_7_9_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_7_9_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_7_9_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_7_9_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_7_9_out_W_noc3_data;
wire tile_7_9_out_N_noc3_valid;
wire tile_7_9_out_S_noc3_valid;
wire tile_7_9_out_E_noc3_valid;
wire tile_7_9_out_W_noc3_valid;
wire tile_7_9_out_N_noc3_yummy;
wire tile_7_9_out_S_noc3_yummy;
wire tile_7_9_out_E_noc3_yummy;
wire tile_7_9_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_8_9_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_8_9_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_8_9_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_8_9_out_W_noc1_data;
wire tile_8_9_out_N_noc1_valid;
wire tile_8_9_out_S_noc1_valid;
wire tile_8_9_out_E_noc1_valid;
wire tile_8_9_out_W_noc1_valid;
wire tile_8_9_out_N_noc1_yummy;
wire tile_8_9_out_S_noc1_yummy;
wire tile_8_9_out_E_noc1_yummy;
wire tile_8_9_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_8_9_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_8_9_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_8_9_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_8_9_out_W_noc2_data;
wire tile_8_9_out_N_noc2_valid;
wire tile_8_9_out_S_noc2_valid;
wire tile_8_9_out_E_noc2_valid;
wire tile_8_9_out_W_noc2_valid;
wire tile_8_9_out_N_noc2_yummy;
wire tile_8_9_out_S_noc2_yummy;
wire tile_8_9_out_E_noc2_yummy;
wire tile_8_9_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_8_9_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_8_9_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_8_9_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_8_9_out_W_noc3_data;
wire tile_8_9_out_N_noc3_valid;
wire tile_8_9_out_S_noc3_valid;
wire tile_8_9_out_E_noc3_valid;
wire tile_8_9_out_W_noc3_valid;
wire tile_8_9_out_N_noc3_yummy;
wire tile_8_9_out_S_noc3_yummy;
wire tile_8_9_out_E_noc3_yummy;
wire tile_8_9_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_9_9_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_9_9_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_9_9_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_9_9_out_W_noc1_data;
wire tile_9_9_out_N_noc1_valid;
wire tile_9_9_out_S_noc1_valid;
wire tile_9_9_out_E_noc1_valid;
wire tile_9_9_out_W_noc1_valid;
wire tile_9_9_out_N_noc1_yummy;
wire tile_9_9_out_S_noc1_yummy;
wire tile_9_9_out_E_noc1_yummy;
wire tile_9_9_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_9_9_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_9_9_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_9_9_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_9_9_out_W_noc2_data;
wire tile_9_9_out_N_noc2_valid;
wire tile_9_9_out_S_noc2_valid;
wire tile_9_9_out_E_noc2_valid;
wire tile_9_9_out_W_noc2_valid;
wire tile_9_9_out_N_noc2_yummy;
wire tile_9_9_out_S_noc2_yummy;
wire tile_9_9_out_E_noc2_yummy;
wire tile_9_9_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_9_9_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_9_9_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_9_9_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_9_9_out_W_noc3_data;
wire tile_9_9_out_N_noc3_valid;
wire tile_9_9_out_S_noc3_valid;
wire tile_9_9_out_E_noc3_valid;
wire tile_9_9_out_W_noc3_valid;
wire tile_9_9_out_N_noc3_yummy;
wire tile_9_9_out_S_noc3_yummy;
wire tile_9_9_out_E_noc3_yummy;
wire tile_9_9_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_10_9_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_10_9_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_10_9_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_10_9_out_W_noc1_data;
wire tile_10_9_out_N_noc1_valid;
wire tile_10_9_out_S_noc1_valid;
wire tile_10_9_out_E_noc1_valid;
wire tile_10_9_out_W_noc1_valid;
wire tile_10_9_out_N_noc1_yummy;
wire tile_10_9_out_S_noc1_yummy;
wire tile_10_9_out_E_noc1_yummy;
wire tile_10_9_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_10_9_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_10_9_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_10_9_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_10_9_out_W_noc2_data;
wire tile_10_9_out_N_noc2_valid;
wire tile_10_9_out_S_noc2_valid;
wire tile_10_9_out_E_noc2_valid;
wire tile_10_9_out_W_noc2_valid;
wire tile_10_9_out_N_noc2_yummy;
wire tile_10_9_out_S_noc2_yummy;
wire tile_10_9_out_E_noc2_yummy;
wire tile_10_9_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_10_9_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_10_9_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_10_9_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_10_9_out_W_noc3_data;
wire tile_10_9_out_N_noc3_valid;
wire tile_10_9_out_S_noc3_valid;
wire tile_10_9_out_E_noc3_valid;
wire tile_10_9_out_W_noc3_valid;
wire tile_10_9_out_N_noc3_yummy;
wire tile_10_9_out_S_noc3_yummy;
wire tile_10_9_out_E_noc3_yummy;
wire tile_10_9_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_11_9_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_11_9_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_11_9_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_11_9_out_W_noc1_data;
wire tile_11_9_out_N_noc1_valid;
wire tile_11_9_out_S_noc1_valid;
wire tile_11_9_out_E_noc1_valid;
wire tile_11_9_out_W_noc1_valid;
wire tile_11_9_out_N_noc1_yummy;
wire tile_11_9_out_S_noc1_yummy;
wire tile_11_9_out_E_noc1_yummy;
wire tile_11_9_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_11_9_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_11_9_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_11_9_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_11_9_out_W_noc2_data;
wire tile_11_9_out_N_noc2_valid;
wire tile_11_9_out_S_noc2_valid;
wire tile_11_9_out_E_noc2_valid;
wire tile_11_9_out_W_noc2_valid;
wire tile_11_9_out_N_noc2_yummy;
wire tile_11_9_out_S_noc2_yummy;
wire tile_11_9_out_E_noc2_yummy;
wire tile_11_9_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_11_9_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_11_9_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_11_9_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_11_9_out_W_noc3_data;
wire tile_11_9_out_N_noc3_valid;
wire tile_11_9_out_S_noc3_valid;
wire tile_11_9_out_E_noc3_valid;
wire tile_11_9_out_W_noc3_valid;
wire tile_11_9_out_N_noc3_yummy;
wire tile_11_9_out_S_noc3_yummy;
wire tile_11_9_out_E_noc3_yummy;
wire tile_11_9_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_12_9_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_12_9_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_12_9_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_12_9_out_W_noc1_data;
wire tile_12_9_out_N_noc1_valid;
wire tile_12_9_out_S_noc1_valid;
wire tile_12_9_out_E_noc1_valid;
wire tile_12_9_out_W_noc1_valid;
wire tile_12_9_out_N_noc1_yummy;
wire tile_12_9_out_S_noc1_yummy;
wire tile_12_9_out_E_noc1_yummy;
wire tile_12_9_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_12_9_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_12_9_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_12_9_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_12_9_out_W_noc2_data;
wire tile_12_9_out_N_noc2_valid;
wire tile_12_9_out_S_noc2_valid;
wire tile_12_9_out_E_noc2_valid;
wire tile_12_9_out_W_noc2_valid;
wire tile_12_9_out_N_noc2_yummy;
wire tile_12_9_out_S_noc2_yummy;
wire tile_12_9_out_E_noc2_yummy;
wire tile_12_9_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_12_9_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_12_9_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_12_9_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_12_9_out_W_noc3_data;
wire tile_12_9_out_N_noc3_valid;
wire tile_12_9_out_S_noc3_valid;
wire tile_12_9_out_E_noc3_valid;
wire tile_12_9_out_W_noc3_valid;
wire tile_12_9_out_N_noc3_yummy;
wire tile_12_9_out_S_noc3_yummy;
wire tile_12_9_out_E_noc3_yummy;
wire tile_12_9_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_13_9_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_13_9_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_13_9_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_13_9_out_W_noc1_data;
wire tile_13_9_out_N_noc1_valid;
wire tile_13_9_out_S_noc1_valid;
wire tile_13_9_out_E_noc1_valid;
wire tile_13_9_out_W_noc1_valid;
wire tile_13_9_out_N_noc1_yummy;
wire tile_13_9_out_S_noc1_yummy;
wire tile_13_9_out_E_noc1_yummy;
wire tile_13_9_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_13_9_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_13_9_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_13_9_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_13_9_out_W_noc2_data;
wire tile_13_9_out_N_noc2_valid;
wire tile_13_9_out_S_noc2_valid;
wire tile_13_9_out_E_noc2_valid;
wire tile_13_9_out_W_noc2_valid;
wire tile_13_9_out_N_noc2_yummy;
wire tile_13_9_out_S_noc2_yummy;
wire tile_13_9_out_E_noc2_yummy;
wire tile_13_9_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_13_9_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_13_9_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_13_9_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_13_9_out_W_noc3_data;
wire tile_13_9_out_N_noc3_valid;
wire tile_13_9_out_S_noc3_valid;
wire tile_13_9_out_E_noc3_valid;
wire tile_13_9_out_W_noc3_valid;
wire tile_13_9_out_N_noc3_yummy;
wire tile_13_9_out_S_noc3_yummy;
wire tile_13_9_out_E_noc3_yummy;
wire tile_13_9_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_14_9_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_14_9_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_14_9_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_14_9_out_W_noc1_data;
wire tile_14_9_out_N_noc1_valid;
wire tile_14_9_out_S_noc1_valid;
wire tile_14_9_out_E_noc1_valid;
wire tile_14_9_out_W_noc1_valid;
wire tile_14_9_out_N_noc1_yummy;
wire tile_14_9_out_S_noc1_yummy;
wire tile_14_9_out_E_noc1_yummy;
wire tile_14_9_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_14_9_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_14_9_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_14_9_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_14_9_out_W_noc2_data;
wire tile_14_9_out_N_noc2_valid;
wire tile_14_9_out_S_noc2_valid;
wire tile_14_9_out_E_noc2_valid;
wire tile_14_9_out_W_noc2_valid;
wire tile_14_9_out_N_noc2_yummy;
wire tile_14_9_out_S_noc2_yummy;
wire tile_14_9_out_E_noc2_yummy;
wire tile_14_9_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_14_9_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_14_9_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_14_9_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_14_9_out_W_noc3_data;
wire tile_14_9_out_N_noc3_valid;
wire tile_14_9_out_S_noc3_valid;
wire tile_14_9_out_E_noc3_valid;
wire tile_14_9_out_W_noc3_valid;
wire tile_14_9_out_N_noc3_yummy;
wire tile_14_9_out_S_noc3_yummy;
wire tile_14_9_out_E_noc3_yummy;
wire tile_14_9_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_15_9_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_15_9_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_15_9_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_15_9_out_W_noc1_data;
wire tile_15_9_out_N_noc1_valid;
wire tile_15_9_out_S_noc1_valid;
wire tile_15_9_out_E_noc1_valid;
wire tile_15_9_out_W_noc1_valid;
wire tile_15_9_out_N_noc1_yummy;
wire tile_15_9_out_S_noc1_yummy;
wire tile_15_9_out_E_noc1_yummy;
wire tile_15_9_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_15_9_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_15_9_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_15_9_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_15_9_out_W_noc2_data;
wire tile_15_9_out_N_noc2_valid;
wire tile_15_9_out_S_noc2_valid;
wire tile_15_9_out_E_noc2_valid;
wire tile_15_9_out_W_noc2_valid;
wire tile_15_9_out_N_noc2_yummy;
wire tile_15_9_out_S_noc2_yummy;
wire tile_15_9_out_E_noc2_yummy;
wire tile_15_9_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_15_9_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_15_9_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_15_9_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_15_9_out_W_noc3_data;
wire tile_15_9_out_N_noc3_valid;
wire tile_15_9_out_S_noc3_valid;
wire tile_15_9_out_E_noc3_valid;
wire tile_15_9_out_W_noc3_valid;
wire tile_15_9_out_N_noc3_yummy;
wire tile_15_9_out_S_noc3_yummy;
wire tile_15_9_out_E_noc3_yummy;
wire tile_15_9_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_0_10_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_0_10_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_0_10_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_0_10_out_W_noc1_data;
wire tile_0_10_out_N_noc1_valid;
wire tile_0_10_out_S_noc1_valid;
wire tile_0_10_out_E_noc1_valid;
wire tile_0_10_out_W_noc1_valid;
wire tile_0_10_out_N_noc1_yummy;
wire tile_0_10_out_S_noc1_yummy;
wire tile_0_10_out_E_noc1_yummy;
wire tile_0_10_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_0_10_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_0_10_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_0_10_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_0_10_out_W_noc2_data;
wire tile_0_10_out_N_noc2_valid;
wire tile_0_10_out_S_noc2_valid;
wire tile_0_10_out_E_noc2_valid;
wire tile_0_10_out_W_noc2_valid;
wire tile_0_10_out_N_noc2_yummy;
wire tile_0_10_out_S_noc2_yummy;
wire tile_0_10_out_E_noc2_yummy;
wire tile_0_10_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_0_10_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_0_10_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_0_10_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_0_10_out_W_noc3_data;
wire tile_0_10_out_N_noc3_valid;
wire tile_0_10_out_S_noc3_valid;
wire tile_0_10_out_E_noc3_valid;
wire tile_0_10_out_W_noc3_valid;
wire tile_0_10_out_N_noc3_yummy;
wire tile_0_10_out_S_noc3_yummy;
wire tile_0_10_out_E_noc3_yummy;
wire tile_0_10_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_1_10_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_1_10_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_1_10_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_1_10_out_W_noc1_data;
wire tile_1_10_out_N_noc1_valid;
wire tile_1_10_out_S_noc1_valid;
wire tile_1_10_out_E_noc1_valid;
wire tile_1_10_out_W_noc1_valid;
wire tile_1_10_out_N_noc1_yummy;
wire tile_1_10_out_S_noc1_yummy;
wire tile_1_10_out_E_noc1_yummy;
wire tile_1_10_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_1_10_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_1_10_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_1_10_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_1_10_out_W_noc2_data;
wire tile_1_10_out_N_noc2_valid;
wire tile_1_10_out_S_noc2_valid;
wire tile_1_10_out_E_noc2_valid;
wire tile_1_10_out_W_noc2_valid;
wire tile_1_10_out_N_noc2_yummy;
wire tile_1_10_out_S_noc2_yummy;
wire tile_1_10_out_E_noc2_yummy;
wire tile_1_10_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_1_10_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_1_10_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_1_10_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_1_10_out_W_noc3_data;
wire tile_1_10_out_N_noc3_valid;
wire tile_1_10_out_S_noc3_valid;
wire tile_1_10_out_E_noc3_valid;
wire tile_1_10_out_W_noc3_valid;
wire tile_1_10_out_N_noc3_yummy;
wire tile_1_10_out_S_noc3_yummy;
wire tile_1_10_out_E_noc3_yummy;
wire tile_1_10_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_2_10_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_2_10_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_2_10_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_2_10_out_W_noc1_data;
wire tile_2_10_out_N_noc1_valid;
wire tile_2_10_out_S_noc1_valid;
wire tile_2_10_out_E_noc1_valid;
wire tile_2_10_out_W_noc1_valid;
wire tile_2_10_out_N_noc1_yummy;
wire tile_2_10_out_S_noc1_yummy;
wire tile_2_10_out_E_noc1_yummy;
wire tile_2_10_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_2_10_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_2_10_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_2_10_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_2_10_out_W_noc2_data;
wire tile_2_10_out_N_noc2_valid;
wire tile_2_10_out_S_noc2_valid;
wire tile_2_10_out_E_noc2_valid;
wire tile_2_10_out_W_noc2_valid;
wire tile_2_10_out_N_noc2_yummy;
wire tile_2_10_out_S_noc2_yummy;
wire tile_2_10_out_E_noc2_yummy;
wire tile_2_10_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_2_10_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_2_10_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_2_10_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_2_10_out_W_noc3_data;
wire tile_2_10_out_N_noc3_valid;
wire tile_2_10_out_S_noc3_valid;
wire tile_2_10_out_E_noc3_valid;
wire tile_2_10_out_W_noc3_valid;
wire tile_2_10_out_N_noc3_yummy;
wire tile_2_10_out_S_noc3_yummy;
wire tile_2_10_out_E_noc3_yummy;
wire tile_2_10_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_3_10_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_3_10_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_3_10_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_3_10_out_W_noc1_data;
wire tile_3_10_out_N_noc1_valid;
wire tile_3_10_out_S_noc1_valid;
wire tile_3_10_out_E_noc1_valid;
wire tile_3_10_out_W_noc1_valid;
wire tile_3_10_out_N_noc1_yummy;
wire tile_3_10_out_S_noc1_yummy;
wire tile_3_10_out_E_noc1_yummy;
wire tile_3_10_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_3_10_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_3_10_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_3_10_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_3_10_out_W_noc2_data;
wire tile_3_10_out_N_noc2_valid;
wire tile_3_10_out_S_noc2_valid;
wire tile_3_10_out_E_noc2_valid;
wire tile_3_10_out_W_noc2_valid;
wire tile_3_10_out_N_noc2_yummy;
wire tile_3_10_out_S_noc2_yummy;
wire tile_3_10_out_E_noc2_yummy;
wire tile_3_10_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_3_10_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_3_10_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_3_10_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_3_10_out_W_noc3_data;
wire tile_3_10_out_N_noc3_valid;
wire tile_3_10_out_S_noc3_valid;
wire tile_3_10_out_E_noc3_valid;
wire tile_3_10_out_W_noc3_valid;
wire tile_3_10_out_N_noc3_yummy;
wire tile_3_10_out_S_noc3_yummy;
wire tile_3_10_out_E_noc3_yummy;
wire tile_3_10_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_4_10_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_4_10_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_4_10_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_4_10_out_W_noc1_data;
wire tile_4_10_out_N_noc1_valid;
wire tile_4_10_out_S_noc1_valid;
wire tile_4_10_out_E_noc1_valid;
wire tile_4_10_out_W_noc1_valid;
wire tile_4_10_out_N_noc1_yummy;
wire tile_4_10_out_S_noc1_yummy;
wire tile_4_10_out_E_noc1_yummy;
wire tile_4_10_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_4_10_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_4_10_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_4_10_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_4_10_out_W_noc2_data;
wire tile_4_10_out_N_noc2_valid;
wire tile_4_10_out_S_noc2_valid;
wire tile_4_10_out_E_noc2_valid;
wire tile_4_10_out_W_noc2_valid;
wire tile_4_10_out_N_noc2_yummy;
wire tile_4_10_out_S_noc2_yummy;
wire tile_4_10_out_E_noc2_yummy;
wire tile_4_10_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_4_10_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_4_10_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_4_10_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_4_10_out_W_noc3_data;
wire tile_4_10_out_N_noc3_valid;
wire tile_4_10_out_S_noc3_valid;
wire tile_4_10_out_E_noc3_valid;
wire tile_4_10_out_W_noc3_valid;
wire tile_4_10_out_N_noc3_yummy;
wire tile_4_10_out_S_noc3_yummy;
wire tile_4_10_out_E_noc3_yummy;
wire tile_4_10_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_5_10_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_5_10_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_5_10_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_5_10_out_W_noc1_data;
wire tile_5_10_out_N_noc1_valid;
wire tile_5_10_out_S_noc1_valid;
wire tile_5_10_out_E_noc1_valid;
wire tile_5_10_out_W_noc1_valid;
wire tile_5_10_out_N_noc1_yummy;
wire tile_5_10_out_S_noc1_yummy;
wire tile_5_10_out_E_noc1_yummy;
wire tile_5_10_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_5_10_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_5_10_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_5_10_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_5_10_out_W_noc2_data;
wire tile_5_10_out_N_noc2_valid;
wire tile_5_10_out_S_noc2_valid;
wire tile_5_10_out_E_noc2_valid;
wire tile_5_10_out_W_noc2_valid;
wire tile_5_10_out_N_noc2_yummy;
wire tile_5_10_out_S_noc2_yummy;
wire tile_5_10_out_E_noc2_yummy;
wire tile_5_10_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_5_10_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_5_10_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_5_10_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_5_10_out_W_noc3_data;
wire tile_5_10_out_N_noc3_valid;
wire tile_5_10_out_S_noc3_valid;
wire tile_5_10_out_E_noc3_valid;
wire tile_5_10_out_W_noc3_valid;
wire tile_5_10_out_N_noc3_yummy;
wire tile_5_10_out_S_noc3_yummy;
wire tile_5_10_out_E_noc3_yummy;
wire tile_5_10_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_6_10_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_6_10_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_6_10_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_6_10_out_W_noc1_data;
wire tile_6_10_out_N_noc1_valid;
wire tile_6_10_out_S_noc1_valid;
wire tile_6_10_out_E_noc1_valid;
wire tile_6_10_out_W_noc1_valid;
wire tile_6_10_out_N_noc1_yummy;
wire tile_6_10_out_S_noc1_yummy;
wire tile_6_10_out_E_noc1_yummy;
wire tile_6_10_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_6_10_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_6_10_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_6_10_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_6_10_out_W_noc2_data;
wire tile_6_10_out_N_noc2_valid;
wire tile_6_10_out_S_noc2_valid;
wire tile_6_10_out_E_noc2_valid;
wire tile_6_10_out_W_noc2_valid;
wire tile_6_10_out_N_noc2_yummy;
wire tile_6_10_out_S_noc2_yummy;
wire tile_6_10_out_E_noc2_yummy;
wire tile_6_10_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_6_10_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_6_10_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_6_10_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_6_10_out_W_noc3_data;
wire tile_6_10_out_N_noc3_valid;
wire tile_6_10_out_S_noc3_valid;
wire tile_6_10_out_E_noc3_valid;
wire tile_6_10_out_W_noc3_valid;
wire tile_6_10_out_N_noc3_yummy;
wire tile_6_10_out_S_noc3_yummy;
wire tile_6_10_out_E_noc3_yummy;
wire tile_6_10_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_7_10_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_7_10_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_7_10_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_7_10_out_W_noc1_data;
wire tile_7_10_out_N_noc1_valid;
wire tile_7_10_out_S_noc1_valid;
wire tile_7_10_out_E_noc1_valid;
wire tile_7_10_out_W_noc1_valid;
wire tile_7_10_out_N_noc1_yummy;
wire tile_7_10_out_S_noc1_yummy;
wire tile_7_10_out_E_noc1_yummy;
wire tile_7_10_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_7_10_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_7_10_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_7_10_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_7_10_out_W_noc2_data;
wire tile_7_10_out_N_noc2_valid;
wire tile_7_10_out_S_noc2_valid;
wire tile_7_10_out_E_noc2_valid;
wire tile_7_10_out_W_noc2_valid;
wire tile_7_10_out_N_noc2_yummy;
wire tile_7_10_out_S_noc2_yummy;
wire tile_7_10_out_E_noc2_yummy;
wire tile_7_10_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_7_10_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_7_10_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_7_10_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_7_10_out_W_noc3_data;
wire tile_7_10_out_N_noc3_valid;
wire tile_7_10_out_S_noc3_valid;
wire tile_7_10_out_E_noc3_valid;
wire tile_7_10_out_W_noc3_valid;
wire tile_7_10_out_N_noc3_yummy;
wire tile_7_10_out_S_noc3_yummy;
wire tile_7_10_out_E_noc3_yummy;
wire tile_7_10_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_8_10_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_8_10_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_8_10_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_8_10_out_W_noc1_data;
wire tile_8_10_out_N_noc1_valid;
wire tile_8_10_out_S_noc1_valid;
wire tile_8_10_out_E_noc1_valid;
wire tile_8_10_out_W_noc1_valid;
wire tile_8_10_out_N_noc1_yummy;
wire tile_8_10_out_S_noc1_yummy;
wire tile_8_10_out_E_noc1_yummy;
wire tile_8_10_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_8_10_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_8_10_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_8_10_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_8_10_out_W_noc2_data;
wire tile_8_10_out_N_noc2_valid;
wire tile_8_10_out_S_noc2_valid;
wire tile_8_10_out_E_noc2_valid;
wire tile_8_10_out_W_noc2_valid;
wire tile_8_10_out_N_noc2_yummy;
wire tile_8_10_out_S_noc2_yummy;
wire tile_8_10_out_E_noc2_yummy;
wire tile_8_10_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_8_10_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_8_10_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_8_10_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_8_10_out_W_noc3_data;
wire tile_8_10_out_N_noc3_valid;
wire tile_8_10_out_S_noc3_valid;
wire tile_8_10_out_E_noc3_valid;
wire tile_8_10_out_W_noc3_valid;
wire tile_8_10_out_N_noc3_yummy;
wire tile_8_10_out_S_noc3_yummy;
wire tile_8_10_out_E_noc3_yummy;
wire tile_8_10_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_9_10_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_9_10_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_9_10_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_9_10_out_W_noc1_data;
wire tile_9_10_out_N_noc1_valid;
wire tile_9_10_out_S_noc1_valid;
wire tile_9_10_out_E_noc1_valid;
wire tile_9_10_out_W_noc1_valid;
wire tile_9_10_out_N_noc1_yummy;
wire tile_9_10_out_S_noc1_yummy;
wire tile_9_10_out_E_noc1_yummy;
wire tile_9_10_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_9_10_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_9_10_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_9_10_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_9_10_out_W_noc2_data;
wire tile_9_10_out_N_noc2_valid;
wire tile_9_10_out_S_noc2_valid;
wire tile_9_10_out_E_noc2_valid;
wire tile_9_10_out_W_noc2_valid;
wire tile_9_10_out_N_noc2_yummy;
wire tile_9_10_out_S_noc2_yummy;
wire tile_9_10_out_E_noc2_yummy;
wire tile_9_10_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_9_10_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_9_10_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_9_10_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_9_10_out_W_noc3_data;
wire tile_9_10_out_N_noc3_valid;
wire tile_9_10_out_S_noc3_valid;
wire tile_9_10_out_E_noc3_valid;
wire tile_9_10_out_W_noc3_valid;
wire tile_9_10_out_N_noc3_yummy;
wire tile_9_10_out_S_noc3_yummy;
wire tile_9_10_out_E_noc3_yummy;
wire tile_9_10_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_10_10_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_10_10_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_10_10_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_10_10_out_W_noc1_data;
wire tile_10_10_out_N_noc1_valid;
wire tile_10_10_out_S_noc1_valid;
wire tile_10_10_out_E_noc1_valid;
wire tile_10_10_out_W_noc1_valid;
wire tile_10_10_out_N_noc1_yummy;
wire tile_10_10_out_S_noc1_yummy;
wire tile_10_10_out_E_noc1_yummy;
wire tile_10_10_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_10_10_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_10_10_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_10_10_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_10_10_out_W_noc2_data;
wire tile_10_10_out_N_noc2_valid;
wire tile_10_10_out_S_noc2_valid;
wire tile_10_10_out_E_noc2_valid;
wire tile_10_10_out_W_noc2_valid;
wire tile_10_10_out_N_noc2_yummy;
wire tile_10_10_out_S_noc2_yummy;
wire tile_10_10_out_E_noc2_yummy;
wire tile_10_10_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_10_10_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_10_10_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_10_10_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_10_10_out_W_noc3_data;
wire tile_10_10_out_N_noc3_valid;
wire tile_10_10_out_S_noc3_valid;
wire tile_10_10_out_E_noc3_valid;
wire tile_10_10_out_W_noc3_valid;
wire tile_10_10_out_N_noc3_yummy;
wire tile_10_10_out_S_noc3_yummy;
wire tile_10_10_out_E_noc3_yummy;
wire tile_10_10_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_11_10_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_11_10_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_11_10_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_11_10_out_W_noc1_data;
wire tile_11_10_out_N_noc1_valid;
wire tile_11_10_out_S_noc1_valid;
wire tile_11_10_out_E_noc1_valid;
wire tile_11_10_out_W_noc1_valid;
wire tile_11_10_out_N_noc1_yummy;
wire tile_11_10_out_S_noc1_yummy;
wire tile_11_10_out_E_noc1_yummy;
wire tile_11_10_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_11_10_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_11_10_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_11_10_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_11_10_out_W_noc2_data;
wire tile_11_10_out_N_noc2_valid;
wire tile_11_10_out_S_noc2_valid;
wire tile_11_10_out_E_noc2_valid;
wire tile_11_10_out_W_noc2_valid;
wire tile_11_10_out_N_noc2_yummy;
wire tile_11_10_out_S_noc2_yummy;
wire tile_11_10_out_E_noc2_yummy;
wire tile_11_10_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_11_10_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_11_10_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_11_10_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_11_10_out_W_noc3_data;
wire tile_11_10_out_N_noc3_valid;
wire tile_11_10_out_S_noc3_valid;
wire tile_11_10_out_E_noc3_valid;
wire tile_11_10_out_W_noc3_valid;
wire tile_11_10_out_N_noc3_yummy;
wire tile_11_10_out_S_noc3_yummy;
wire tile_11_10_out_E_noc3_yummy;
wire tile_11_10_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_12_10_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_12_10_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_12_10_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_12_10_out_W_noc1_data;
wire tile_12_10_out_N_noc1_valid;
wire tile_12_10_out_S_noc1_valid;
wire tile_12_10_out_E_noc1_valid;
wire tile_12_10_out_W_noc1_valid;
wire tile_12_10_out_N_noc1_yummy;
wire tile_12_10_out_S_noc1_yummy;
wire tile_12_10_out_E_noc1_yummy;
wire tile_12_10_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_12_10_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_12_10_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_12_10_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_12_10_out_W_noc2_data;
wire tile_12_10_out_N_noc2_valid;
wire tile_12_10_out_S_noc2_valid;
wire tile_12_10_out_E_noc2_valid;
wire tile_12_10_out_W_noc2_valid;
wire tile_12_10_out_N_noc2_yummy;
wire tile_12_10_out_S_noc2_yummy;
wire tile_12_10_out_E_noc2_yummy;
wire tile_12_10_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_12_10_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_12_10_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_12_10_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_12_10_out_W_noc3_data;
wire tile_12_10_out_N_noc3_valid;
wire tile_12_10_out_S_noc3_valid;
wire tile_12_10_out_E_noc3_valid;
wire tile_12_10_out_W_noc3_valid;
wire tile_12_10_out_N_noc3_yummy;
wire tile_12_10_out_S_noc3_yummy;
wire tile_12_10_out_E_noc3_yummy;
wire tile_12_10_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_13_10_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_13_10_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_13_10_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_13_10_out_W_noc1_data;
wire tile_13_10_out_N_noc1_valid;
wire tile_13_10_out_S_noc1_valid;
wire tile_13_10_out_E_noc1_valid;
wire tile_13_10_out_W_noc1_valid;
wire tile_13_10_out_N_noc1_yummy;
wire tile_13_10_out_S_noc1_yummy;
wire tile_13_10_out_E_noc1_yummy;
wire tile_13_10_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_13_10_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_13_10_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_13_10_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_13_10_out_W_noc2_data;
wire tile_13_10_out_N_noc2_valid;
wire tile_13_10_out_S_noc2_valid;
wire tile_13_10_out_E_noc2_valid;
wire tile_13_10_out_W_noc2_valid;
wire tile_13_10_out_N_noc2_yummy;
wire tile_13_10_out_S_noc2_yummy;
wire tile_13_10_out_E_noc2_yummy;
wire tile_13_10_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_13_10_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_13_10_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_13_10_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_13_10_out_W_noc3_data;
wire tile_13_10_out_N_noc3_valid;
wire tile_13_10_out_S_noc3_valid;
wire tile_13_10_out_E_noc3_valid;
wire tile_13_10_out_W_noc3_valid;
wire tile_13_10_out_N_noc3_yummy;
wire tile_13_10_out_S_noc3_yummy;
wire tile_13_10_out_E_noc3_yummy;
wire tile_13_10_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_14_10_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_14_10_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_14_10_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_14_10_out_W_noc1_data;
wire tile_14_10_out_N_noc1_valid;
wire tile_14_10_out_S_noc1_valid;
wire tile_14_10_out_E_noc1_valid;
wire tile_14_10_out_W_noc1_valid;
wire tile_14_10_out_N_noc1_yummy;
wire tile_14_10_out_S_noc1_yummy;
wire tile_14_10_out_E_noc1_yummy;
wire tile_14_10_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_14_10_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_14_10_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_14_10_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_14_10_out_W_noc2_data;
wire tile_14_10_out_N_noc2_valid;
wire tile_14_10_out_S_noc2_valid;
wire tile_14_10_out_E_noc2_valid;
wire tile_14_10_out_W_noc2_valid;
wire tile_14_10_out_N_noc2_yummy;
wire tile_14_10_out_S_noc2_yummy;
wire tile_14_10_out_E_noc2_yummy;
wire tile_14_10_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_14_10_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_14_10_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_14_10_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_14_10_out_W_noc3_data;
wire tile_14_10_out_N_noc3_valid;
wire tile_14_10_out_S_noc3_valid;
wire tile_14_10_out_E_noc3_valid;
wire tile_14_10_out_W_noc3_valid;
wire tile_14_10_out_N_noc3_yummy;
wire tile_14_10_out_S_noc3_yummy;
wire tile_14_10_out_E_noc3_yummy;
wire tile_14_10_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_15_10_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_15_10_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_15_10_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_15_10_out_W_noc1_data;
wire tile_15_10_out_N_noc1_valid;
wire tile_15_10_out_S_noc1_valid;
wire tile_15_10_out_E_noc1_valid;
wire tile_15_10_out_W_noc1_valid;
wire tile_15_10_out_N_noc1_yummy;
wire tile_15_10_out_S_noc1_yummy;
wire tile_15_10_out_E_noc1_yummy;
wire tile_15_10_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_15_10_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_15_10_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_15_10_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_15_10_out_W_noc2_data;
wire tile_15_10_out_N_noc2_valid;
wire tile_15_10_out_S_noc2_valid;
wire tile_15_10_out_E_noc2_valid;
wire tile_15_10_out_W_noc2_valid;
wire tile_15_10_out_N_noc2_yummy;
wire tile_15_10_out_S_noc2_yummy;
wire tile_15_10_out_E_noc2_yummy;
wire tile_15_10_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_15_10_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_15_10_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_15_10_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_15_10_out_W_noc3_data;
wire tile_15_10_out_N_noc3_valid;
wire tile_15_10_out_S_noc3_valid;
wire tile_15_10_out_E_noc3_valid;
wire tile_15_10_out_W_noc3_valid;
wire tile_15_10_out_N_noc3_yummy;
wire tile_15_10_out_S_noc3_yummy;
wire tile_15_10_out_E_noc3_yummy;
wire tile_15_10_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_0_11_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_0_11_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_0_11_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_0_11_out_W_noc1_data;
wire tile_0_11_out_N_noc1_valid;
wire tile_0_11_out_S_noc1_valid;
wire tile_0_11_out_E_noc1_valid;
wire tile_0_11_out_W_noc1_valid;
wire tile_0_11_out_N_noc1_yummy;
wire tile_0_11_out_S_noc1_yummy;
wire tile_0_11_out_E_noc1_yummy;
wire tile_0_11_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_0_11_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_0_11_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_0_11_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_0_11_out_W_noc2_data;
wire tile_0_11_out_N_noc2_valid;
wire tile_0_11_out_S_noc2_valid;
wire tile_0_11_out_E_noc2_valid;
wire tile_0_11_out_W_noc2_valid;
wire tile_0_11_out_N_noc2_yummy;
wire tile_0_11_out_S_noc2_yummy;
wire tile_0_11_out_E_noc2_yummy;
wire tile_0_11_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_0_11_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_0_11_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_0_11_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_0_11_out_W_noc3_data;
wire tile_0_11_out_N_noc3_valid;
wire tile_0_11_out_S_noc3_valid;
wire tile_0_11_out_E_noc3_valid;
wire tile_0_11_out_W_noc3_valid;
wire tile_0_11_out_N_noc3_yummy;
wire tile_0_11_out_S_noc3_yummy;
wire tile_0_11_out_E_noc3_yummy;
wire tile_0_11_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_1_11_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_1_11_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_1_11_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_1_11_out_W_noc1_data;
wire tile_1_11_out_N_noc1_valid;
wire tile_1_11_out_S_noc1_valid;
wire tile_1_11_out_E_noc1_valid;
wire tile_1_11_out_W_noc1_valid;
wire tile_1_11_out_N_noc1_yummy;
wire tile_1_11_out_S_noc1_yummy;
wire tile_1_11_out_E_noc1_yummy;
wire tile_1_11_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_1_11_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_1_11_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_1_11_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_1_11_out_W_noc2_data;
wire tile_1_11_out_N_noc2_valid;
wire tile_1_11_out_S_noc2_valid;
wire tile_1_11_out_E_noc2_valid;
wire tile_1_11_out_W_noc2_valid;
wire tile_1_11_out_N_noc2_yummy;
wire tile_1_11_out_S_noc2_yummy;
wire tile_1_11_out_E_noc2_yummy;
wire tile_1_11_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_1_11_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_1_11_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_1_11_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_1_11_out_W_noc3_data;
wire tile_1_11_out_N_noc3_valid;
wire tile_1_11_out_S_noc3_valid;
wire tile_1_11_out_E_noc3_valid;
wire tile_1_11_out_W_noc3_valid;
wire tile_1_11_out_N_noc3_yummy;
wire tile_1_11_out_S_noc3_yummy;
wire tile_1_11_out_E_noc3_yummy;
wire tile_1_11_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_2_11_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_2_11_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_2_11_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_2_11_out_W_noc1_data;
wire tile_2_11_out_N_noc1_valid;
wire tile_2_11_out_S_noc1_valid;
wire tile_2_11_out_E_noc1_valid;
wire tile_2_11_out_W_noc1_valid;
wire tile_2_11_out_N_noc1_yummy;
wire tile_2_11_out_S_noc1_yummy;
wire tile_2_11_out_E_noc1_yummy;
wire tile_2_11_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_2_11_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_2_11_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_2_11_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_2_11_out_W_noc2_data;
wire tile_2_11_out_N_noc2_valid;
wire tile_2_11_out_S_noc2_valid;
wire tile_2_11_out_E_noc2_valid;
wire tile_2_11_out_W_noc2_valid;
wire tile_2_11_out_N_noc2_yummy;
wire tile_2_11_out_S_noc2_yummy;
wire tile_2_11_out_E_noc2_yummy;
wire tile_2_11_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_2_11_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_2_11_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_2_11_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_2_11_out_W_noc3_data;
wire tile_2_11_out_N_noc3_valid;
wire tile_2_11_out_S_noc3_valid;
wire tile_2_11_out_E_noc3_valid;
wire tile_2_11_out_W_noc3_valid;
wire tile_2_11_out_N_noc3_yummy;
wire tile_2_11_out_S_noc3_yummy;
wire tile_2_11_out_E_noc3_yummy;
wire tile_2_11_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_3_11_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_3_11_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_3_11_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_3_11_out_W_noc1_data;
wire tile_3_11_out_N_noc1_valid;
wire tile_3_11_out_S_noc1_valid;
wire tile_3_11_out_E_noc1_valid;
wire tile_3_11_out_W_noc1_valid;
wire tile_3_11_out_N_noc1_yummy;
wire tile_3_11_out_S_noc1_yummy;
wire tile_3_11_out_E_noc1_yummy;
wire tile_3_11_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_3_11_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_3_11_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_3_11_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_3_11_out_W_noc2_data;
wire tile_3_11_out_N_noc2_valid;
wire tile_3_11_out_S_noc2_valid;
wire tile_3_11_out_E_noc2_valid;
wire tile_3_11_out_W_noc2_valid;
wire tile_3_11_out_N_noc2_yummy;
wire tile_3_11_out_S_noc2_yummy;
wire tile_3_11_out_E_noc2_yummy;
wire tile_3_11_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_3_11_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_3_11_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_3_11_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_3_11_out_W_noc3_data;
wire tile_3_11_out_N_noc3_valid;
wire tile_3_11_out_S_noc3_valid;
wire tile_3_11_out_E_noc3_valid;
wire tile_3_11_out_W_noc3_valid;
wire tile_3_11_out_N_noc3_yummy;
wire tile_3_11_out_S_noc3_yummy;
wire tile_3_11_out_E_noc3_yummy;
wire tile_3_11_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_4_11_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_4_11_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_4_11_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_4_11_out_W_noc1_data;
wire tile_4_11_out_N_noc1_valid;
wire tile_4_11_out_S_noc1_valid;
wire tile_4_11_out_E_noc1_valid;
wire tile_4_11_out_W_noc1_valid;
wire tile_4_11_out_N_noc1_yummy;
wire tile_4_11_out_S_noc1_yummy;
wire tile_4_11_out_E_noc1_yummy;
wire tile_4_11_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_4_11_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_4_11_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_4_11_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_4_11_out_W_noc2_data;
wire tile_4_11_out_N_noc2_valid;
wire tile_4_11_out_S_noc2_valid;
wire tile_4_11_out_E_noc2_valid;
wire tile_4_11_out_W_noc2_valid;
wire tile_4_11_out_N_noc2_yummy;
wire tile_4_11_out_S_noc2_yummy;
wire tile_4_11_out_E_noc2_yummy;
wire tile_4_11_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_4_11_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_4_11_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_4_11_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_4_11_out_W_noc3_data;
wire tile_4_11_out_N_noc3_valid;
wire tile_4_11_out_S_noc3_valid;
wire tile_4_11_out_E_noc3_valid;
wire tile_4_11_out_W_noc3_valid;
wire tile_4_11_out_N_noc3_yummy;
wire tile_4_11_out_S_noc3_yummy;
wire tile_4_11_out_E_noc3_yummy;
wire tile_4_11_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_5_11_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_5_11_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_5_11_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_5_11_out_W_noc1_data;
wire tile_5_11_out_N_noc1_valid;
wire tile_5_11_out_S_noc1_valid;
wire tile_5_11_out_E_noc1_valid;
wire tile_5_11_out_W_noc1_valid;
wire tile_5_11_out_N_noc1_yummy;
wire tile_5_11_out_S_noc1_yummy;
wire tile_5_11_out_E_noc1_yummy;
wire tile_5_11_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_5_11_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_5_11_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_5_11_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_5_11_out_W_noc2_data;
wire tile_5_11_out_N_noc2_valid;
wire tile_5_11_out_S_noc2_valid;
wire tile_5_11_out_E_noc2_valid;
wire tile_5_11_out_W_noc2_valid;
wire tile_5_11_out_N_noc2_yummy;
wire tile_5_11_out_S_noc2_yummy;
wire tile_5_11_out_E_noc2_yummy;
wire tile_5_11_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_5_11_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_5_11_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_5_11_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_5_11_out_W_noc3_data;
wire tile_5_11_out_N_noc3_valid;
wire tile_5_11_out_S_noc3_valid;
wire tile_5_11_out_E_noc3_valid;
wire tile_5_11_out_W_noc3_valid;
wire tile_5_11_out_N_noc3_yummy;
wire tile_5_11_out_S_noc3_yummy;
wire tile_5_11_out_E_noc3_yummy;
wire tile_5_11_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_6_11_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_6_11_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_6_11_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_6_11_out_W_noc1_data;
wire tile_6_11_out_N_noc1_valid;
wire tile_6_11_out_S_noc1_valid;
wire tile_6_11_out_E_noc1_valid;
wire tile_6_11_out_W_noc1_valid;
wire tile_6_11_out_N_noc1_yummy;
wire tile_6_11_out_S_noc1_yummy;
wire tile_6_11_out_E_noc1_yummy;
wire tile_6_11_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_6_11_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_6_11_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_6_11_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_6_11_out_W_noc2_data;
wire tile_6_11_out_N_noc2_valid;
wire tile_6_11_out_S_noc2_valid;
wire tile_6_11_out_E_noc2_valid;
wire tile_6_11_out_W_noc2_valid;
wire tile_6_11_out_N_noc2_yummy;
wire tile_6_11_out_S_noc2_yummy;
wire tile_6_11_out_E_noc2_yummy;
wire tile_6_11_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_6_11_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_6_11_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_6_11_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_6_11_out_W_noc3_data;
wire tile_6_11_out_N_noc3_valid;
wire tile_6_11_out_S_noc3_valid;
wire tile_6_11_out_E_noc3_valid;
wire tile_6_11_out_W_noc3_valid;
wire tile_6_11_out_N_noc3_yummy;
wire tile_6_11_out_S_noc3_yummy;
wire tile_6_11_out_E_noc3_yummy;
wire tile_6_11_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_7_11_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_7_11_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_7_11_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_7_11_out_W_noc1_data;
wire tile_7_11_out_N_noc1_valid;
wire tile_7_11_out_S_noc1_valid;
wire tile_7_11_out_E_noc1_valid;
wire tile_7_11_out_W_noc1_valid;
wire tile_7_11_out_N_noc1_yummy;
wire tile_7_11_out_S_noc1_yummy;
wire tile_7_11_out_E_noc1_yummy;
wire tile_7_11_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_7_11_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_7_11_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_7_11_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_7_11_out_W_noc2_data;
wire tile_7_11_out_N_noc2_valid;
wire tile_7_11_out_S_noc2_valid;
wire tile_7_11_out_E_noc2_valid;
wire tile_7_11_out_W_noc2_valid;
wire tile_7_11_out_N_noc2_yummy;
wire tile_7_11_out_S_noc2_yummy;
wire tile_7_11_out_E_noc2_yummy;
wire tile_7_11_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_7_11_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_7_11_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_7_11_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_7_11_out_W_noc3_data;
wire tile_7_11_out_N_noc3_valid;
wire tile_7_11_out_S_noc3_valid;
wire tile_7_11_out_E_noc3_valid;
wire tile_7_11_out_W_noc3_valid;
wire tile_7_11_out_N_noc3_yummy;
wire tile_7_11_out_S_noc3_yummy;
wire tile_7_11_out_E_noc3_yummy;
wire tile_7_11_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_8_11_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_8_11_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_8_11_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_8_11_out_W_noc1_data;
wire tile_8_11_out_N_noc1_valid;
wire tile_8_11_out_S_noc1_valid;
wire tile_8_11_out_E_noc1_valid;
wire tile_8_11_out_W_noc1_valid;
wire tile_8_11_out_N_noc1_yummy;
wire tile_8_11_out_S_noc1_yummy;
wire tile_8_11_out_E_noc1_yummy;
wire tile_8_11_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_8_11_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_8_11_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_8_11_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_8_11_out_W_noc2_data;
wire tile_8_11_out_N_noc2_valid;
wire tile_8_11_out_S_noc2_valid;
wire tile_8_11_out_E_noc2_valid;
wire tile_8_11_out_W_noc2_valid;
wire tile_8_11_out_N_noc2_yummy;
wire tile_8_11_out_S_noc2_yummy;
wire tile_8_11_out_E_noc2_yummy;
wire tile_8_11_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_8_11_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_8_11_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_8_11_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_8_11_out_W_noc3_data;
wire tile_8_11_out_N_noc3_valid;
wire tile_8_11_out_S_noc3_valid;
wire tile_8_11_out_E_noc3_valid;
wire tile_8_11_out_W_noc3_valid;
wire tile_8_11_out_N_noc3_yummy;
wire tile_8_11_out_S_noc3_yummy;
wire tile_8_11_out_E_noc3_yummy;
wire tile_8_11_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_9_11_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_9_11_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_9_11_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_9_11_out_W_noc1_data;
wire tile_9_11_out_N_noc1_valid;
wire tile_9_11_out_S_noc1_valid;
wire tile_9_11_out_E_noc1_valid;
wire tile_9_11_out_W_noc1_valid;
wire tile_9_11_out_N_noc1_yummy;
wire tile_9_11_out_S_noc1_yummy;
wire tile_9_11_out_E_noc1_yummy;
wire tile_9_11_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_9_11_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_9_11_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_9_11_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_9_11_out_W_noc2_data;
wire tile_9_11_out_N_noc2_valid;
wire tile_9_11_out_S_noc2_valid;
wire tile_9_11_out_E_noc2_valid;
wire tile_9_11_out_W_noc2_valid;
wire tile_9_11_out_N_noc2_yummy;
wire tile_9_11_out_S_noc2_yummy;
wire tile_9_11_out_E_noc2_yummy;
wire tile_9_11_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_9_11_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_9_11_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_9_11_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_9_11_out_W_noc3_data;
wire tile_9_11_out_N_noc3_valid;
wire tile_9_11_out_S_noc3_valid;
wire tile_9_11_out_E_noc3_valid;
wire tile_9_11_out_W_noc3_valid;
wire tile_9_11_out_N_noc3_yummy;
wire tile_9_11_out_S_noc3_yummy;
wire tile_9_11_out_E_noc3_yummy;
wire tile_9_11_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_10_11_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_10_11_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_10_11_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_10_11_out_W_noc1_data;
wire tile_10_11_out_N_noc1_valid;
wire tile_10_11_out_S_noc1_valid;
wire tile_10_11_out_E_noc1_valid;
wire tile_10_11_out_W_noc1_valid;
wire tile_10_11_out_N_noc1_yummy;
wire tile_10_11_out_S_noc1_yummy;
wire tile_10_11_out_E_noc1_yummy;
wire tile_10_11_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_10_11_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_10_11_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_10_11_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_10_11_out_W_noc2_data;
wire tile_10_11_out_N_noc2_valid;
wire tile_10_11_out_S_noc2_valid;
wire tile_10_11_out_E_noc2_valid;
wire tile_10_11_out_W_noc2_valid;
wire tile_10_11_out_N_noc2_yummy;
wire tile_10_11_out_S_noc2_yummy;
wire tile_10_11_out_E_noc2_yummy;
wire tile_10_11_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_10_11_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_10_11_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_10_11_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_10_11_out_W_noc3_data;
wire tile_10_11_out_N_noc3_valid;
wire tile_10_11_out_S_noc3_valid;
wire tile_10_11_out_E_noc3_valid;
wire tile_10_11_out_W_noc3_valid;
wire tile_10_11_out_N_noc3_yummy;
wire tile_10_11_out_S_noc3_yummy;
wire tile_10_11_out_E_noc3_yummy;
wire tile_10_11_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_11_11_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_11_11_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_11_11_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_11_11_out_W_noc1_data;
wire tile_11_11_out_N_noc1_valid;
wire tile_11_11_out_S_noc1_valid;
wire tile_11_11_out_E_noc1_valid;
wire tile_11_11_out_W_noc1_valid;
wire tile_11_11_out_N_noc1_yummy;
wire tile_11_11_out_S_noc1_yummy;
wire tile_11_11_out_E_noc1_yummy;
wire tile_11_11_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_11_11_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_11_11_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_11_11_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_11_11_out_W_noc2_data;
wire tile_11_11_out_N_noc2_valid;
wire tile_11_11_out_S_noc2_valid;
wire tile_11_11_out_E_noc2_valid;
wire tile_11_11_out_W_noc2_valid;
wire tile_11_11_out_N_noc2_yummy;
wire tile_11_11_out_S_noc2_yummy;
wire tile_11_11_out_E_noc2_yummy;
wire tile_11_11_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_11_11_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_11_11_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_11_11_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_11_11_out_W_noc3_data;
wire tile_11_11_out_N_noc3_valid;
wire tile_11_11_out_S_noc3_valid;
wire tile_11_11_out_E_noc3_valid;
wire tile_11_11_out_W_noc3_valid;
wire tile_11_11_out_N_noc3_yummy;
wire tile_11_11_out_S_noc3_yummy;
wire tile_11_11_out_E_noc3_yummy;
wire tile_11_11_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_12_11_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_12_11_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_12_11_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_12_11_out_W_noc1_data;
wire tile_12_11_out_N_noc1_valid;
wire tile_12_11_out_S_noc1_valid;
wire tile_12_11_out_E_noc1_valid;
wire tile_12_11_out_W_noc1_valid;
wire tile_12_11_out_N_noc1_yummy;
wire tile_12_11_out_S_noc1_yummy;
wire tile_12_11_out_E_noc1_yummy;
wire tile_12_11_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_12_11_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_12_11_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_12_11_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_12_11_out_W_noc2_data;
wire tile_12_11_out_N_noc2_valid;
wire tile_12_11_out_S_noc2_valid;
wire tile_12_11_out_E_noc2_valid;
wire tile_12_11_out_W_noc2_valid;
wire tile_12_11_out_N_noc2_yummy;
wire tile_12_11_out_S_noc2_yummy;
wire tile_12_11_out_E_noc2_yummy;
wire tile_12_11_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_12_11_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_12_11_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_12_11_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_12_11_out_W_noc3_data;
wire tile_12_11_out_N_noc3_valid;
wire tile_12_11_out_S_noc3_valid;
wire tile_12_11_out_E_noc3_valid;
wire tile_12_11_out_W_noc3_valid;
wire tile_12_11_out_N_noc3_yummy;
wire tile_12_11_out_S_noc3_yummy;
wire tile_12_11_out_E_noc3_yummy;
wire tile_12_11_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_13_11_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_13_11_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_13_11_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_13_11_out_W_noc1_data;
wire tile_13_11_out_N_noc1_valid;
wire tile_13_11_out_S_noc1_valid;
wire tile_13_11_out_E_noc1_valid;
wire tile_13_11_out_W_noc1_valid;
wire tile_13_11_out_N_noc1_yummy;
wire tile_13_11_out_S_noc1_yummy;
wire tile_13_11_out_E_noc1_yummy;
wire tile_13_11_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_13_11_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_13_11_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_13_11_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_13_11_out_W_noc2_data;
wire tile_13_11_out_N_noc2_valid;
wire tile_13_11_out_S_noc2_valid;
wire tile_13_11_out_E_noc2_valid;
wire tile_13_11_out_W_noc2_valid;
wire tile_13_11_out_N_noc2_yummy;
wire tile_13_11_out_S_noc2_yummy;
wire tile_13_11_out_E_noc2_yummy;
wire tile_13_11_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_13_11_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_13_11_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_13_11_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_13_11_out_W_noc3_data;
wire tile_13_11_out_N_noc3_valid;
wire tile_13_11_out_S_noc3_valid;
wire tile_13_11_out_E_noc3_valid;
wire tile_13_11_out_W_noc3_valid;
wire tile_13_11_out_N_noc3_yummy;
wire tile_13_11_out_S_noc3_yummy;
wire tile_13_11_out_E_noc3_yummy;
wire tile_13_11_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_14_11_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_14_11_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_14_11_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_14_11_out_W_noc1_data;
wire tile_14_11_out_N_noc1_valid;
wire tile_14_11_out_S_noc1_valid;
wire tile_14_11_out_E_noc1_valid;
wire tile_14_11_out_W_noc1_valid;
wire tile_14_11_out_N_noc1_yummy;
wire tile_14_11_out_S_noc1_yummy;
wire tile_14_11_out_E_noc1_yummy;
wire tile_14_11_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_14_11_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_14_11_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_14_11_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_14_11_out_W_noc2_data;
wire tile_14_11_out_N_noc2_valid;
wire tile_14_11_out_S_noc2_valid;
wire tile_14_11_out_E_noc2_valid;
wire tile_14_11_out_W_noc2_valid;
wire tile_14_11_out_N_noc2_yummy;
wire tile_14_11_out_S_noc2_yummy;
wire tile_14_11_out_E_noc2_yummy;
wire tile_14_11_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_14_11_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_14_11_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_14_11_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_14_11_out_W_noc3_data;
wire tile_14_11_out_N_noc3_valid;
wire tile_14_11_out_S_noc3_valid;
wire tile_14_11_out_E_noc3_valid;
wire tile_14_11_out_W_noc3_valid;
wire tile_14_11_out_N_noc3_yummy;
wire tile_14_11_out_S_noc3_yummy;
wire tile_14_11_out_E_noc3_yummy;
wire tile_14_11_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_15_11_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_15_11_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_15_11_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_15_11_out_W_noc1_data;
wire tile_15_11_out_N_noc1_valid;
wire tile_15_11_out_S_noc1_valid;
wire tile_15_11_out_E_noc1_valid;
wire tile_15_11_out_W_noc1_valid;
wire tile_15_11_out_N_noc1_yummy;
wire tile_15_11_out_S_noc1_yummy;
wire tile_15_11_out_E_noc1_yummy;
wire tile_15_11_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_15_11_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_15_11_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_15_11_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_15_11_out_W_noc2_data;
wire tile_15_11_out_N_noc2_valid;
wire tile_15_11_out_S_noc2_valid;
wire tile_15_11_out_E_noc2_valid;
wire tile_15_11_out_W_noc2_valid;
wire tile_15_11_out_N_noc2_yummy;
wire tile_15_11_out_S_noc2_yummy;
wire tile_15_11_out_E_noc2_yummy;
wire tile_15_11_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_15_11_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_15_11_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_15_11_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_15_11_out_W_noc3_data;
wire tile_15_11_out_N_noc3_valid;
wire tile_15_11_out_S_noc3_valid;
wire tile_15_11_out_E_noc3_valid;
wire tile_15_11_out_W_noc3_valid;
wire tile_15_11_out_N_noc3_yummy;
wire tile_15_11_out_S_noc3_yummy;
wire tile_15_11_out_E_noc3_yummy;
wire tile_15_11_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_0_12_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_0_12_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_0_12_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_0_12_out_W_noc1_data;
wire tile_0_12_out_N_noc1_valid;
wire tile_0_12_out_S_noc1_valid;
wire tile_0_12_out_E_noc1_valid;
wire tile_0_12_out_W_noc1_valid;
wire tile_0_12_out_N_noc1_yummy;
wire tile_0_12_out_S_noc1_yummy;
wire tile_0_12_out_E_noc1_yummy;
wire tile_0_12_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_0_12_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_0_12_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_0_12_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_0_12_out_W_noc2_data;
wire tile_0_12_out_N_noc2_valid;
wire tile_0_12_out_S_noc2_valid;
wire tile_0_12_out_E_noc2_valid;
wire tile_0_12_out_W_noc2_valid;
wire tile_0_12_out_N_noc2_yummy;
wire tile_0_12_out_S_noc2_yummy;
wire tile_0_12_out_E_noc2_yummy;
wire tile_0_12_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_0_12_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_0_12_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_0_12_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_0_12_out_W_noc3_data;
wire tile_0_12_out_N_noc3_valid;
wire tile_0_12_out_S_noc3_valid;
wire tile_0_12_out_E_noc3_valid;
wire tile_0_12_out_W_noc3_valid;
wire tile_0_12_out_N_noc3_yummy;
wire tile_0_12_out_S_noc3_yummy;
wire tile_0_12_out_E_noc3_yummy;
wire tile_0_12_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_1_12_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_1_12_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_1_12_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_1_12_out_W_noc1_data;
wire tile_1_12_out_N_noc1_valid;
wire tile_1_12_out_S_noc1_valid;
wire tile_1_12_out_E_noc1_valid;
wire tile_1_12_out_W_noc1_valid;
wire tile_1_12_out_N_noc1_yummy;
wire tile_1_12_out_S_noc1_yummy;
wire tile_1_12_out_E_noc1_yummy;
wire tile_1_12_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_1_12_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_1_12_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_1_12_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_1_12_out_W_noc2_data;
wire tile_1_12_out_N_noc2_valid;
wire tile_1_12_out_S_noc2_valid;
wire tile_1_12_out_E_noc2_valid;
wire tile_1_12_out_W_noc2_valid;
wire tile_1_12_out_N_noc2_yummy;
wire tile_1_12_out_S_noc2_yummy;
wire tile_1_12_out_E_noc2_yummy;
wire tile_1_12_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_1_12_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_1_12_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_1_12_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_1_12_out_W_noc3_data;
wire tile_1_12_out_N_noc3_valid;
wire tile_1_12_out_S_noc3_valid;
wire tile_1_12_out_E_noc3_valid;
wire tile_1_12_out_W_noc3_valid;
wire tile_1_12_out_N_noc3_yummy;
wire tile_1_12_out_S_noc3_yummy;
wire tile_1_12_out_E_noc3_yummy;
wire tile_1_12_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_2_12_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_2_12_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_2_12_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_2_12_out_W_noc1_data;
wire tile_2_12_out_N_noc1_valid;
wire tile_2_12_out_S_noc1_valid;
wire tile_2_12_out_E_noc1_valid;
wire tile_2_12_out_W_noc1_valid;
wire tile_2_12_out_N_noc1_yummy;
wire tile_2_12_out_S_noc1_yummy;
wire tile_2_12_out_E_noc1_yummy;
wire tile_2_12_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_2_12_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_2_12_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_2_12_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_2_12_out_W_noc2_data;
wire tile_2_12_out_N_noc2_valid;
wire tile_2_12_out_S_noc2_valid;
wire tile_2_12_out_E_noc2_valid;
wire tile_2_12_out_W_noc2_valid;
wire tile_2_12_out_N_noc2_yummy;
wire tile_2_12_out_S_noc2_yummy;
wire tile_2_12_out_E_noc2_yummy;
wire tile_2_12_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_2_12_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_2_12_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_2_12_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_2_12_out_W_noc3_data;
wire tile_2_12_out_N_noc3_valid;
wire tile_2_12_out_S_noc3_valid;
wire tile_2_12_out_E_noc3_valid;
wire tile_2_12_out_W_noc3_valid;
wire tile_2_12_out_N_noc3_yummy;
wire tile_2_12_out_S_noc3_yummy;
wire tile_2_12_out_E_noc3_yummy;
wire tile_2_12_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_3_12_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_3_12_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_3_12_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_3_12_out_W_noc1_data;
wire tile_3_12_out_N_noc1_valid;
wire tile_3_12_out_S_noc1_valid;
wire tile_3_12_out_E_noc1_valid;
wire tile_3_12_out_W_noc1_valid;
wire tile_3_12_out_N_noc1_yummy;
wire tile_3_12_out_S_noc1_yummy;
wire tile_3_12_out_E_noc1_yummy;
wire tile_3_12_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_3_12_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_3_12_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_3_12_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_3_12_out_W_noc2_data;
wire tile_3_12_out_N_noc2_valid;
wire tile_3_12_out_S_noc2_valid;
wire tile_3_12_out_E_noc2_valid;
wire tile_3_12_out_W_noc2_valid;
wire tile_3_12_out_N_noc2_yummy;
wire tile_3_12_out_S_noc2_yummy;
wire tile_3_12_out_E_noc2_yummy;
wire tile_3_12_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_3_12_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_3_12_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_3_12_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_3_12_out_W_noc3_data;
wire tile_3_12_out_N_noc3_valid;
wire tile_3_12_out_S_noc3_valid;
wire tile_3_12_out_E_noc3_valid;
wire tile_3_12_out_W_noc3_valid;
wire tile_3_12_out_N_noc3_yummy;
wire tile_3_12_out_S_noc3_yummy;
wire tile_3_12_out_E_noc3_yummy;
wire tile_3_12_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_4_12_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_4_12_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_4_12_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_4_12_out_W_noc1_data;
wire tile_4_12_out_N_noc1_valid;
wire tile_4_12_out_S_noc1_valid;
wire tile_4_12_out_E_noc1_valid;
wire tile_4_12_out_W_noc1_valid;
wire tile_4_12_out_N_noc1_yummy;
wire tile_4_12_out_S_noc1_yummy;
wire tile_4_12_out_E_noc1_yummy;
wire tile_4_12_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_4_12_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_4_12_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_4_12_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_4_12_out_W_noc2_data;
wire tile_4_12_out_N_noc2_valid;
wire tile_4_12_out_S_noc2_valid;
wire tile_4_12_out_E_noc2_valid;
wire tile_4_12_out_W_noc2_valid;
wire tile_4_12_out_N_noc2_yummy;
wire tile_4_12_out_S_noc2_yummy;
wire tile_4_12_out_E_noc2_yummy;
wire tile_4_12_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_4_12_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_4_12_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_4_12_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_4_12_out_W_noc3_data;
wire tile_4_12_out_N_noc3_valid;
wire tile_4_12_out_S_noc3_valid;
wire tile_4_12_out_E_noc3_valid;
wire tile_4_12_out_W_noc3_valid;
wire tile_4_12_out_N_noc3_yummy;
wire tile_4_12_out_S_noc3_yummy;
wire tile_4_12_out_E_noc3_yummy;
wire tile_4_12_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_5_12_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_5_12_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_5_12_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_5_12_out_W_noc1_data;
wire tile_5_12_out_N_noc1_valid;
wire tile_5_12_out_S_noc1_valid;
wire tile_5_12_out_E_noc1_valid;
wire tile_5_12_out_W_noc1_valid;
wire tile_5_12_out_N_noc1_yummy;
wire tile_5_12_out_S_noc1_yummy;
wire tile_5_12_out_E_noc1_yummy;
wire tile_5_12_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_5_12_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_5_12_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_5_12_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_5_12_out_W_noc2_data;
wire tile_5_12_out_N_noc2_valid;
wire tile_5_12_out_S_noc2_valid;
wire tile_5_12_out_E_noc2_valid;
wire tile_5_12_out_W_noc2_valid;
wire tile_5_12_out_N_noc2_yummy;
wire tile_5_12_out_S_noc2_yummy;
wire tile_5_12_out_E_noc2_yummy;
wire tile_5_12_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_5_12_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_5_12_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_5_12_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_5_12_out_W_noc3_data;
wire tile_5_12_out_N_noc3_valid;
wire tile_5_12_out_S_noc3_valid;
wire tile_5_12_out_E_noc3_valid;
wire tile_5_12_out_W_noc3_valid;
wire tile_5_12_out_N_noc3_yummy;
wire tile_5_12_out_S_noc3_yummy;
wire tile_5_12_out_E_noc3_yummy;
wire tile_5_12_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_6_12_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_6_12_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_6_12_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_6_12_out_W_noc1_data;
wire tile_6_12_out_N_noc1_valid;
wire tile_6_12_out_S_noc1_valid;
wire tile_6_12_out_E_noc1_valid;
wire tile_6_12_out_W_noc1_valid;
wire tile_6_12_out_N_noc1_yummy;
wire tile_6_12_out_S_noc1_yummy;
wire tile_6_12_out_E_noc1_yummy;
wire tile_6_12_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_6_12_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_6_12_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_6_12_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_6_12_out_W_noc2_data;
wire tile_6_12_out_N_noc2_valid;
wire tile_6_12_out_S_noc2_valid;
wire tile_6_12_out_E_noc2_valid;
wire tile_6_12_out_W_noc2_valid;
wire tile_6_12_out_N_noc2_yummy;
wire tile_6_12_out_S_noc2_yummy;
wire tile_6_12_out_E_noc2_yummy;
wire tile_6_12_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_6_12_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_6_12_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_6_12_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_6_12_out_W_noc3_data;
wire tile_6_12_out_N_noc3_valid;
wire tile_6_12_out_S_noc3_valid;
wire tile_6_12_out_E_noc3_valid;
wire tile_6_12_out_W_noc3_valid;
wire tile_6_12_out_N_noc3_yummy;
wire tile_6_12_out_S_noc3_yummy;
wire tile_6_12_out_E_noc3_yummy;
wire tile_6_12_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_7_12_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_7_12_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_7_12_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_7_12_out_W_noc1_data;
wire tile_7_12_out_N_noc1_valid;
wire tile_7_12_out_S_noc1_valid;
wire tile_7_12_out_E_noc1_valid;
wire tile_7_12_out_W_noc1_valid;
wire tile_7_12_out_N_noc1_yummy;
wire tile_7_12_out_S_noc1_yummy;
wire tile_7_12_out_E_noc1_yummy;
wire tile_7_12_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_7_12_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_7_12_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_7_12_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_7_12_out_W_noc2_data;
wire tile_7_12_out_N_noc2_valid;
wire tile_7_12_out_S_noc2_valid;
wire tile_7_12_out_E_noc2_valid;
wire tile_7_12_out_W_noc2_valid;
wire tile_7_12_out_N_noc2_yummy;
wire tile_7_12_out_S_noc2_yummy;
wire tile_7_12_out_E_noc2_yummy;
wire tile_7_12_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_7_12_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_7_12_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_7_12_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_7_12_out_W_noc3_data;
wire tile_7_12_out_N_noc3_valid;
wire tile_7_12_out_S_noc3_valid;
wire tile_7_12_out_E_noc3_valid;
wire tile_7_12_out_W_noc3_valid;
wire tile_7_12_out_N_noc3_yummy;
wire tile_7_12_out_S_noc3_yummy;
wire tile_7_12_out_E_noc3_yummy;
wire tile_7_12_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_8_12_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_8_12_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_8_12_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_8_12_out_W_noc1_data;
wire tile_8_12_out_N_noc1_valid;
wire tile_8_12_out_S_noc1_valid;
wire tile_8_12_out_E_noc1_valid;
wire tile_8_12_out_W_noc1_valid;
wire tile_8_12_out_N_noc1_yummy;
wire tile_8_12_out_S_noc1_yummy;
wire tile_8_12_out_E_noc1_yummy;
wire tile_8_12_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_8_12_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_8_12_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_8_12_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_8_12_out_W_noc2_data;
wire tile_8_12_out_N_noc2_valid;
wire tile_8_12_out_S_noc2_valid;
wire tile_8_12_out_E_noc2_valid;
wire tile_8_12_out_W_noc2_valid;
wire tile_8_12_out_N_noc2_yummy;
wire tile_8_12_out_S_noc2_yummy;
wire tile_8_12_out_E_noc2_yummy;
wire tile_8_12_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_8_12_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_8_12_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_8_12_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_8_12_out_W_noc3_data;
wire tile_8_12_out_N_noc3_valid;
wire tile_8_12_out_S_noc3_valid;
wire tile_8_12_out_E_noc3_valid;
wire tile_8_12_out_W_noc3_valid;
wire tile_8_12_out_N_noc3_yummy;
wire tile_8_12_out_S_noc3_yummy;
wire tile_8_12_out_E_noc3_yummy;
wire tile_8_12_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_9_12_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_9_12_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_9_12_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_9_12_out_W_noc1_data;
wire tile_9_12_out_N_noc1_valid;
wire tile_9_12_out_S_noc1_valid;
wire tile_9_12_out_E_noc1_valid;
wire tile_9_12_out_W_noc1_valid;
wire tile_9_12_out_N_noc1_yummy;
wire tile_9_12_out_S_noc1_yummy;
wire tile_9_12_out_E_noc1_yummy;
wire tile_9_12_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_9_12_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_9_12_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_9_12_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_9_12_out_W_noc2_data;
wire tile_9_12_out_N_noc2_valid;
wire tile_9_12_out_S_noc2_valid;
wire tile_9_12_out_E_noc2_valid;
wire tile_9_12_out_W_noc2_valid;
wire tile_9_12_out_N_noc2_yummy;
wire tile_9_12_out_S_noc2_yummy;
wire tile_9_12_out_E_noc2_yummy;
wire tile_9_12_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_9_12_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_9_12_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_9_12_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_9_12_out_W_noc3_data;
wire tile_9_12_out_N_noc3_valid;
wire tile_9_12_out_S_noc3_valid;
wire tile_9_12_out_E_noc3_valid;
wire tile_9_12_out_W_noc3_valid;
wire tile_9_12_out_N_noc3_yummy;
wire tile_9_12_out_S_noc3_yummy;
wire tile_9_12_out_E_noc3_yummy;
wire tile_9_12_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_10_12_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_10_12_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_10_12_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_10_12_out_W_noc1_data;
wire tile_10_12_out_N_noc1_valid;
wire tile_10_12_out_S_noc1_valid;
wire tile_10_12_out_E_noc1_valid;
wire tile_10_12_out_W_noc1_valid;
wire tile_10_12_out_N_noc1_yummy;
wire tile_10_12_out_S_noc1_yummy;
wire tile_10_12_out_E_noc1_yummy;
wire tile_10_12_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_10_12_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_10_12_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_10_12_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_10_12_out_W_noc2_data;
wire tile_10_12_out_N_noc2_valid;
wire tile_10_12_out_S_noc2_valid;
wire tile_10_12_out_E_noc2_valid;
wire tile_10_12_out_W_noc2_valid;
wire tile_10_12_out_N_noc2_yummy;
wire tile_10_12_out_S_noc2_yummy;
wire tile_10_12_out_E_noc2_yummy;
wire tile_10_12_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_10_12_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_10_12_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_10_12_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_10_12_out_W_noc3_data;
wire tile_10_12_out_N_noc3_valid;
wire tile_10_12_out_S_noc3_valid;
wire tile_10_12_out_E_noc3_valid;
wire tile_10_12_out_W_noc3_valid;
wire tile_10_12_out_N_noc3_yummy;
wire tile_10_12_out_S_noc3_yummy;
wire tile_10_12_out_E_noc3_yummy;
wire tile_10_12_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_11_12_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_11_12_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_11_12_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_11_12_out_W_noc1_data;
wire tile_11_12_out_N_noc1_valid;
wire tile_11_12_out_S_noc1_valid;
wire tile_11_12_out_E_noc1_valid;
wire tile_11_12_out_W_noc1_valid;
wire tile_11_12_out_N_noc1_yummy;
wire tile_11_12_out_S_noc1_yummy;
wire tile_11_12_out_E_noc1_yummy;
wire tile_11_12_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_11_12_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_11_12_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_11_12_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_11_12_out_W_noc2_data;
wire tile_11_12_out_N_noc2_valid;
wire tile_11_12_out_S_noc2_valid;
wire tile_11_12_out_E_noc2_valid;
wire tile_11_12_out_W_noc2_valid;
wire tile_11_12_out_N_noc2_yummy;
wire tile_11_12_out_S_noc2_yummy;
wire tile_11_12_out_E_noc2_yummy;
wire tile_11_12_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_11_12_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_11_12_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_11_12_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_11_12_out_W_noc3_data;
wire tile_11_12_out_N_noc3_valid;
wire tile_11_12_out_S_noc3_valid;
wire tile_11_12_out_E_noc3_valid;
wire tile_11_12_out_W_noc3_valid;
wire tile_11_12_out_N_noc3_yummy;
wire tile_11_12_out_S_noc3_yummy;
wire tile_11_12_out_E_noc3_yummy;
wire tile_11_12_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_12_12_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_12_12_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_12_12_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_12_12_out_W_noc1_data;
wire tile_12_12_out_N_noc1_valid;
wire tile_12_12_out_S_noc1_valid;
wire tile_12_12_out_E_noc1_valid;
wire tile_12_12_out_W_noc1_valid;
wire tile_12_12_out_N_noc1_yummy;
wire tile_12_12_out_S_noc1_yummy;
wire tile_12_12_out_E_noc1_yummy;
wire tile_12_12_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_12_12_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_12_12_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_12_12_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_12_12_out_W_noc2_data;
wire tile_12_12_out_N_noc2_valid;
wire tile_12_12_out_S_noc2_valid;
wire tile_12_12_out_E_noc2_valid;
wire tile_12_12_out_W_noc2_valid;
wire tile_12_12_out_N_noc2_yummy;
wire tile_12_12_out_S_noc2_yummy;
wire tile_12_12_out_E_noc2_yummy;
wire tile_12_12_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_12_12_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_12_12_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_12_12_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_12_12_out_W_noc3_data;
wire tile_12_12_out_N_noc3_valid;
wire tile_12_12_out_S_noc3_valid;
wire tile_12_12_out_E_noc3_valid;
wire tile_12_12_out_W_noc3_valid;
wire tile_12_12_out_N_noc3_yummy;
wire tile_12_12_out_S_noc3_yummy;
wire tile_12_12_out_E_noc3_yummy;
wire tile_12_12_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_13_12_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_13_12_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_13_12_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_13_12_out_W_noc1_data;
wire tile_13_12_out_N_noc1_valid;
wire tile_13_12_out_S_noc1_valid;
wire tile_13_12_out_E_noc1_valid;
wire tile_13_12_out_W_noc1_valid;
wire tile_13_12_out_N_noc1_yummy;
wire tile_13_12_out_S_noc1_yummy;
wire tile_13_12_out_E_noc1_yummy;
wire tile_13_12_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_13_12_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_13_12_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_13_12_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_13_12_out_W_noc2_data;
wire tile_13_12_out_N_noc2_valid;
wire tile_13_12_out_S_noc2_valid;
wire tile_13_12_out_E_noc2_valid;
wire tile_13_12_out_W_noc2_valid;
wire tile_13_12_out_N_noc2_yummy;
wire tile_13_12_out_S_noc2_yummy;
wire tile_13_12_out_E_noc2_yummy;
wire tile_13_12_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_13_12_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_13_12_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_13_12_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_13_12_out_W_noc3_data;
wire tile_13_12_out_N_noc3_valid;
wire tile_13_12_out_S_noc3_valid;
wire tile_13_12_out_E_noc3_valid;
wire tile_13_12_out_W_noc3_valid;
wire tile_13_12_out_N_noc3_yummy;
wire tile_13_12_out_S_noc3_yummy;
wire tile_13_12_out_E_noc3_yummy;
wire tile_13_12_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_14_12_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_14_12_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_14_12_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_14_12_out_W_noc1_data;
wire tile_14_12_out_N_noc1_valid;
wire tile_14_12_out_S_noc1_valid;
wire tile_14_12_out_E_noc1_valid;
wire tile_14_12_out_W_noc1_valid;
wire tile_14_12_out_N_noc1_yummy;
wire tile_14_12_out_S_noc1_yummy;
wire tile_14_12_out_E_noc1_yummy;
wire tile_14_12_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_14_12_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_14_12_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_14_12_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_14_12_out_W_noc2_data;
wire tile_14_12_out_N_noc2_valid;
wire tile_14_12_out_S_noc2_valid;
wire tile_14_12_out_E_noc2_valid;
wire tile_14_12_out_W_noc2_valid;
wire tile_14_12_out_N_noc2_yummy;
wire tile_14_12_out_S_noc2_yummy;
wire tile_14_12_out_E_noc2_yummy;
wire tile_14_12_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_14_12_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_14_12_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_14_12_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_14_12_out_W_noc3_data;
wire tile_14_12_out_N_noc3_valid;
wire tile_14_12_out_S_noc3_valid;
wire tile_14_12_out_E_noc3_valid;
wire tile_14_12_out_W_noc3_valid;
wire tile_14_12_out_N_noc3_yummy;
wire tile_14_12_out_S_noc3_yummy;
wire tile_14_12_out_E_noc3_yummy;
wire tile_14_12_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_15_12_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_15_12_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_15_12_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_15_12_out_W_noc1_data;
wire tile_15_12_out_N_noc1_valid;
wire tile_15_12_out_S_noc1_valid;
wire tile_15_12_out_E_noc1_valid;
wire tile_15_12_out_W_noc1_valid;
wire tile_15_12_out_N_noc1_yummy;
wire tile_15_12_out_S_noc1_yummy;
wire tile_15_12_out_E_noc1_yummy;
wire tile_15_12_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_15_12_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_15_12_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_15_12_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_15_12_out_W_noc2_data;
wire tile_15_12_out_N_noc2_valid;
wire tile_15_12_out_S_noc2_valid;
wire tile_15_12_out_E_noc2_valid;
wire tile_15_12_out_W_noc2_valid;
wire tile_15_12_out_N_noc2_yummy;
wire tile_15_12_out_S_noc2_yummy;
wire tile_15_12_out_E_noc2_yummy;
wire tile_15_12_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_15_12_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_15_12_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_15_12_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_15_12_out_W_noc3_data;
wire tile_15_12_out_N_noc3_valid;
wire tile_15_12_out_S_noc3_valid;
wire tile_15_12_out_E_noc3_valid;
wire tile_15_12_out_W_noc3_valid;
wire tile_15_12_out_N_noc3_yummy;
wire tile_15_12_out_S_noc3_yummy;
wire tile_15_12_out_E_noc3_yummy;
wire tile_15_12_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_0_13_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_0_13_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_0_13_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_0_13_out_W_noc1_data;
wire tile_0_13_out_N_noc1_valid;
wire tile_0_13_out_S_noc1_valid;
wire tile_0_13_out_E_noc1_valid;
wire tile_0_13_out_W_noc1_valid;
wire tile_0_13_out_N_noc1_yummy;
wire tile_0_13_out_S_noc1_yummy;
wire tile_0_13_out_E_noc1_yummy;
wire tile_0_13_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_0_13_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_0_13_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_0_13_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_0_13_out_W_noc2_data;
wire tile_0_13_out_N_noc2_valid;
wire tile_0_13_out_S_noc2_valid;
wire tile_0_13_out_E_noc2_valid;
wire tile_0_13_out_W_noc2_valid;
wire tile_0_13_out_N_noc2_yummy;
wire tile_0_13_out_S_noc2_yummy;
wire tile_0_13_out_E_noc2_yummy;
wire tile_0_13_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_0_13_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_0_13_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_0_13_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_0_13_out_W_noc3_data;
wire tile_0_13_out_N_noc3_valid;
wire tile_0_13_out_S_noc3_valid;
wire tile_0_13_out_E_noc3_valid;
wire tile_0_13_out_W_noc3_valid;
wire tile_0_13_out_N_noc3_yummy;
wire tile_0_13_out_S_noc3_yummy;
wire tile_0_13_out_E_noc3_yummy;
wire tile_0_13_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_1_13_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_1_13_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_1_13_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_1_13_out_W_noc1_data;
wire tile_1_13_out_N_noc1_valid;
wire tile_1_13_out_S_noc1_valid;
wire tile_1_13_out_E_noc1_valid;
wire tile_1_13_out_W_noc1_valid;
wire tile_1_13_out_N_noc1_yummy;
wire tile_1_13_out_S_noc1_yummy;
wire tile_1_13_out_E_noc1_yummy;
wire tile_1_13_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_1_13_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_1_13_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_1_13_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_1_13_out_W_noc2_data;
wire tile_1_13_out_N_noc2_valid;
wire tile_1_13_out_S_noc2_valid;
wire tile_1_13_out_E_noc2_valid;
wire tile_1_13_out_W_noc2_valid;
wire tile_1_13_out_N_noc2_yummy;
wire tile_1_13_out_S_noc2_yummy;
wire tile_1_13_out_E_noc2_yummy;
wire tile_1_13_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_1_13_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_1_13_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_1_13_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_1_13_out_W_noc3_data;
wire tile_1_13_out_N_noc3_valid;
wire tile_1_13_out_S_noc3_valid;
wire tile_1_13_out_E_noc3_valid;
wire tile_1_13_out_W_noc3_valid;
wire tile_1_13_out_N_noc3_yummy;
wire tile_1_13_out_S_noc3_yummy;
wire tile_1_13_out_E_noc3_yummy;
wire tile_1_13_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_2_13_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_2_13_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_2_13_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_2_13_out_W_noc1_data;
wire tile_2_13_out_N_noc1_valid;
wire tile_2_13_out_S_noc1_valid;
wire tile_2_13_out_E_noc1_valid;
wire tile_2_13_out_W_noc1_valid;
wire tile_2_13_out_N_noc1_yummy;
wire tile_2_13_out_S_noc1_yummy;
wire tile_2_13_out_E_noc1_yummy;
wire tile_2_13_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_2_13_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_2_13_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_2_13_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_2_13_out_W_noc2_data;
wire tile_2_13_out_N_noc2_valid;
wire tile_2_13_out_S_noc2_valid;
wire tile_2_13_out_E_noc2_valid;
wire tile_2_13_out_W_noc2_valid;
wire tile_2_13_out_N_noc2_yummy;
wire tile_2_13_out_S_noc2_yummy;
wire tile_2_13_out_E_noc2_yummy;
wire tile_2_13_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_2_13_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_2_13_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_2_13_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_2_13_out_W_noc3_data;
wire tile_2_13_out_N_noc3_valid;
wire tile_2_13_out_S_noc3_valid;
wire tile_2_13_out_E_noc3_valid;
wire tile_2_13_out_W_noc3_valid;
wire tile_2_13_out_N_noc3_yummy;
wire tile_2_13_out_S_noc3_yummy;
wire tile_2_13_out_E_noc3_yummy;
wire tile_2_13_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_3_13_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_3_13_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_3_13_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_3_13_out_W_noc1_data;
wire tile_3_13_out_N_noc1_valid;
wire tile_3_13_out_S_noc1_valid;
wire tile_3_13_out_E_noc1_valid;
wire tile_3_13_out_W_noc1_valid;
wire tile_3_13_out_N_noc1_yummy;
wire tile_3_13_out_S_noc1_yummy;
wire tile_3_13_out_E_noc1_yummy;
wire tile_3_13_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_3_13_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_3_13_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_3_13_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_3_13_out_W_noc2_data;
wire tile_3_13_out_N_noc2_valid;
wire tile_3_13_out_S_noc2_valid;
wire tile_3_13_out_E_noc2_valid;
wire tile_3_13_out_W_noc2_valid;
wire tile_3_13_out_N_noc2_yummy;
wire tile_3_13_out_S_noc2_yummy;
wire tile_3_13_out_E_noc2_yummy;
wire tile_3_13_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_3_13_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_3_13_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_3_13_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_3_13_out_W_noc3_data;
wire tile_3_13_out_N_noc3_valid;
wire tile_3_13_out_S_noc3_valid;
wire tile_3_13_out_E_noc3_valid;
wire tile_3_13_out_W_noc3_valid;
wire tile_3_13_out_N_noc3_yummy;
wire tile_3_13_out_S_noc3_yummy;
wire tile_3_13_out_E_noc3_yummy;
wire tile_3_13_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_4_13_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_4_13_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_4_13_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_4_13_out_W_noc1_data;
wire tile_4_13_out_N_noc1_valid;
wire tile_4_13_out_S_noc1_valid;
wire tile_4_13_out_E_noc1_valid;
wire tile_4_13_out_W_noc1_valid;
wire tile_4_13_out_N_noc1_yummy;
wire tile_4_13_out_S_noc1_yummy;
wire tile_4_13_out_E_noc1_yummy;
wire tile_4_13_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_4_13_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_4_13_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_4_13_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_4_13_out_W_noc2_data;
wire tile_4_13_out_N_noc2_valid;
wire tile_4_13_out_S_noc2_valid;
wire tile_4_13_out_E_noc2_valid;
wire tile_4_13_out_W_noc2_valid;
wire tile_4_13_out_N_noc2_yummy;
wire tile_4_13_out_S_noc2_yummy;
wire tile_4_13_out_E_noc2_yummy;
wire tile_4_13_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_4_13_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_4_13_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_4_13_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_4_13_out_W_noc3_data;
wire tile_4_13_out_N_noc3_valid;
wire tile_4_13_out_S_noc3_valid;
wire tile_4_13_out_E_noc3_valid;
wire tile_4_13_out_W_noc3_valid;
wire tile_4_13_out_N_noc3_yummy;
wire tile_4_13_out_S_noc3_yummy;
wire tile_4_13_out_E_noc3_yummy;
wire tile_4_13_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_5_13_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_5_13_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_5_13_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_5_13_out_W_noc1_data;
wire tile_5_13_out_N_noc1_valid;
wire tile_5_13_out_S_noc1_valid;
wire tile_5_13_out_E_noc1_valid;
wire tile_5_13_out_W_noc1_valid;
wire tile_5_13_out_N_noc1_yummy;
wire tile_5_13_out_S_noc1_yummy;
wire tile_5_13_out_E_noc1_yummy;
wire tile_5_13_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_5_13_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_5_13_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_5_13_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_5_13_out_W_noc2_data;
wire tile_5_13_out_N_noc2_valid;
wire tile_5_13_out_S_noc2_valid;
wire tile_5_13_out_E_noc2_valid;
wire tile_5_13_out_W_noc2_valid;
wire tile_5_13_out_N_noc2_yummy;
wire tile_5_13_out_S_noc2_yummy;
wire tile_5_13_out_E_noc2_yummy;
wire tile_5_13_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_5_13_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_5_13_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_5_13_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_5_13_out_W_noc3_data;
wire tile_5_13_out_N_noc3_valid;
wire tile_5_13_out_S_noc3_valid;
wire tile_5_13_out_E_noc3_valid;
wire tile_5_13_out_W_noc3_valid;
wire tile_5_13_out_N_noc3_yummy;
wire tile_5_13_out_S_noc3_yummy;
wire tile_5_13_out_E_noc3_yummy;
wire tile_5_13_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_6_13_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_6_13_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_6_13_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_6_13_out_W_noc1_data;
wire tile_6_13_out_N_noc1_valid;
wire tile_6_13_out_S_noc1_valid;
wire tile_6_13_out_E_noc1_valid;
wire tile_6_13_out_W_noc1_valid;
wire tile_6_13_out_N_noc1_yummy;
wire tile_6_13_out_S_noc1_yummy;
wire tile_6_13_out_E_noc1_yummy;
wire tile_6_13_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_6_13_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_6_13_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_6_13_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_6_13_out_W_noc2_data;
wire tile_6_13_out_N_noc2_valid;
wire tile_6_13_out_S_noc2_valid;
wire tile_6_13_out_E_noc2_valid;
wire tile_6_13_out_W_noc2_valid;
wire tile_6_13_out_N_noc2_yummy;
wire tile_6_13_out_S_noc2_yummy;
wire tile_6_13_out_E_noc2_yummy;
wire tile_6_13_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_6_13_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_6_13_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_6_13_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_6_13_out_W_noc3_data;
wire tile_6_13_out_N_noc3_valid;
wire tile_6_13_out_S_noc3_valid;
wire tile_6_13_out_E_noc3_valid;
wire tile_6_13_out_W_noc3_valid;
wire tile_6_13_out_N_noc3_yummy;
wire tile_6_13_out_S_noc3_yummy;
wire tile_6_13_out_E_noc3_yummy;
wire tile_6_13_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_7_13_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_7_13_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_7_13_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_7_13_out_W_noc1_data;
wire tile_7_13_out_N_noc1_valid;
wire tile_7_13_out_S_noc1_valid;
wire tile_7_13_out_E_noc1_valid;
wire tile_7_13_out_W_noc1_valid;
wire tile_7_13_out_N_noc1_yummy;
wire tile_7_13_out_S_noc1_yummy;
wire tile_7_13_out_E_noc1_yummy;
wire tile_7_13_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_7_13_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_7_13_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_7_13_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_7_13_out_W_noc2_data;
wire tile_7_13_out_N_noc2_valid;
wire tile_7_13_out_S_noc2_valid;
wire tile_7_13_out_E_noc2_valid;
wire tile_7_13_out_W_noc2_valid;
wire tile_7_13_out_N_noc2_yummy;
wire tile_7_13_out_S_noc2_yummy;
wire tile_7_13_out_E_noc2_yummy;
wire tile_7_13_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_7_13_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_7_13_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_7_13_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_7_13_out_W_noc3_data;
wire tile_7_13_out_N_noc3_valid;
wire tile_7_13_out_S_noc3_valid;
wire tile_7_13_out_E_noc3_valid;
wire tile_7_13_out_W_noc3_valid;
wire tile_7_13_out_N_noc3_yummy;
wire tile_7_13_out_S_noc3_yummy;
wire tile_7_13_out_E_noc3_yummy;
wire tile_7_13_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_8_13_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_8_13_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_8_13_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_8_13_out_W_noc1_data;
wire tile_8_13_out_N_noc1_valid;
wire tile_8_13_out_S_noc1_valid;
wire tile_8_13_out_E_noc1_valid;
wire tile_8_13_out_W_noc1_valid;
wire tile_8_13_out_N_noc1_yummy;
wire tile_8_13_out_S_noc1_yummy;
wire tile_8_13_out_E_noc1_yummy;
wire tile_8_13_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_8_13_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_8_13_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_8_13_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_8_13_out_W_noc2_data;
wire tile_8_13_out_N_noc2_valid;
wire tile_8_13_out_S_noc2_valid;
wire tile_8_13_out_E_noc2_valid;
wire tile_8_13_out_W_noc2_valid;
wire tile_8_13_out_N_noc2_yummy;
wire tile_8_13_out_S_noc2_yummy;
wire tile_8_13_out_E_noc2_yummy;
wire tile_8_13_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_8_13_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_8_13_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_8_13_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_8_13_out_W_noc3_data;
wire tile_8_13_out_N_noc3_valid;
wire tile_8_13_out_S_noc3_valid;
wire tile_8_13_out_E_noc3_valid;
wire tile_8_13_out_W_noc3_valid;
wire tile_8_13_out_N_noc3_yummy;
wire tile_8_13_out_S_noc3_yummy;
wire tile_8_13_out_E_noc3_yummy;
wire tile_8_13_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_9_13_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_9_13_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_9_13_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_9_13_out_W_noc1_data;
wire tile_9_13_out_N_noc1_valid;
wire tile_9_13_out_S_noc1_valid;
wire tile_9_13_out_E_noc1_valid;
wire tile_9_13_out_W_noc1_valid;
wire tile_9_13_out_N_noc1_yummy;
wire tile_9_13_out_S_noc1_yummy;
wire tile_9_13_out_E_noc1_yummy;
wire tile_9_13_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_9_13_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_9_13_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_9_13_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_9_13_out_W_noc2_data;
wire tile_9_13_out_N_noc2_valid;
wire tile_9_13_out_S_noc2_valid;
wire tile_9_13_out_E_noc2_valid;
wire tile_9_13_out_W_noc2_valid;
wire tile_9_13_out_N_noc2_yummy;
wire tile_9_13_out_S_noc2_yummy;
wire tile_9_13_out_E_noc2_yummy;
wire tile_9_13_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_9_13_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_9_13_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_9_13_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_9_13_out_W_noc3_data;
wire tile_9_13_out_N_noc3_valid;
wire tile_9_13_out_S_noc3_valid;
wire tile_9_13_out_E_noc3_valid;
wire tile_9_13_out_W_noc3_valid;
wire tile_9_13_out_N_noc3_yummy;
wire tile_9_13_out_S_noc3_yummy;
wire tile_9_13_out_E_noc3_yummy;
wire tile_9_13_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_10_13_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_10_13_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_10_13_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_10_13_out_W_noc1_data;
wire tile_10_13_out_N_noc1_valid;
wire tile_10_13_out_S_noc1_valid;
wire tile_10_13_out_E_noc1_valid;
wire tile_10_13_out_W_noc1_valid;
wire tile_10_13_out_N_noc1_yummy;
wire tile_10_13_out_S_noc1_yummy;
wire tile_10_13_out_E_noc1_yummy;
wire tile_10_13_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_10_13_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_10_13_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_10_13_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_10_13_out_W_noc2_data;
wire tile_10_13_out_N_noc2_valid;
wire tile_10_13_out_S_noc2_valid;
wire tile_10_13_out_E_noc2_valid;
wire tile_10_13_out_W_noc2_valid;
wire tile_10_13_out_N_noc2_yummy;
wire tile_10_13_out_S_noc2_yummy;
wire tile_10_13_out_E_noc2_yummy;
wire tile_10_13_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_10_13_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_10_13_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_10_13_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_10_13_out_W_noc3_data;
wire tile_10_13_out_N_noc3_valid;
wire tile_10_13_out_S_noc3_valid;
wire tile_10_13_out_E_noc3_valid;
wire tile_10_13_out_W_noc3_valid;
wire tile_10_13_out_N_noc3_yummy;
wire tile_10_13_out_S_noc3_yummy;
wire tile_10_13_out_E_noc3_yummy;
wire tile_10_13_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_11_13_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_11_13_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_11_13_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_11_13_out_W_noc1_data;
wire tile_11_13_out_N_noc1_valid;
wire tile_11_13_out_S_noc1_valid;
wire tile_11_13_out_E_noc1_valid;
wire tile_11_13_out_W_noc1_valid;
wire tile_11_13_out_N_noc1_yummy;
wire tile_11_13_out_S_noc1_yummy;
wire tile_11_13_out_E_noc1_yummy;
wire tile_11_13_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_11_13_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_11_13_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_11_13_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_11_13_out_W_noc2_data;
wire tile_11_13_out_N_noc2_valid;
wire tile_11_13_out_S_noc2_valid;
wire tile_11_13_out_E_noc2_valid;
wire tile_11_13_out_W_noc2_valid;
wire tile_11_13_out_N_noc2_yummy;
wire tile_11_13_out_S_noc2_yummy;
wire tile_11_13_out_E_noc2_yummy;
wire tile_11_13_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_11_13_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_11_13_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_11_13_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_11_13_out_W_noc3_data;
wire tile_11_13_out_N_noc3_valid;
wire tile_11_13_out_S_noc3_valid;
wire tile_11_13_out_E_noc3_valid;
wire tile_11_13_out_W_noc3_valid;
wire tile_11_13_out_N_noc3_yummy;
wire tile_11_13_out_S_noc3_yummy;
wire tile_11_13_out_E_noc3_yummy;
wire tile_11_13_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_12_13_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_12_13_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_12_13_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_12_13_out_W_noc1_data;
wire tile_12_13_out_N_noc1_valid;
wire tile_12_13_out_S_noc1_valid;
wire tile_12_13_out_E_noc1_valid;
wire tile_12_13_out_W_noc1_valid;
wire tile_12_13_out_N_noc1_yummy;
wire tile_12_13_out_S_noc1_yummy;
wire tile_12_13_out_E_noc1_yummy;
wire tile_12_13_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_12_13_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_12_13_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_12_13_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_12_13_out_W_noc2_data;
wire tile_12_13_out_N_noc2_valid;
wire tile_12_13_out_S_noc2_valid;
wire tile_12_13_out_E_noc2_valid;
wire tile_12_13_out_W_noc2_valid;
wire tile_12_13_out_N_noc2_yummy;
wire tile_12_13_out_S_noc2_yummy;
wire tile_12_13_out_E_noc2_yummy;
wire tile_12_13_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_12_13_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_12_13_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_12_13_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_12_13_out_W_noc3_data;
wire tile_12_13_out_N_noc3_valid;
wire tile_12_13_out_S_noc3_valid;
wire tile_12_13_out_E_noc3_valid;
wire tile_12_13_out_W_noc3_valid;
wire tile_12_13_out_N_noc3_yummy;
wire tile_12_13_out_S_noc3_yummy;
wire tile_12_13_out_E_noc3_yummy;
wire tile_12_13_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_13_13_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_13_13_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_13_13_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_13_13_out_W_noc1_data;
wire tile_13_13_out_N_noc1_valid;
wire tile_13_13_out_S_noc1_valid;
wire tile_13_13_out_E_noc1_valid;
wire tile_13_13_out_W_noc1_valid;
wire tile_13_13_out_N_noc1_yummy;
wire tile_13_13_out_S_noc1_yummy;
wire tile_13_13_out_E_noc1_yummy;
wire tile_13_13_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_13_13_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_13_13_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_13_13_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_13_13_out_W_noc2_data;
wire tile_13_13_out_N_noc2_valid;
wire tile_13_13_out_S_noc2_valid;
wire tile_13_13_out_E_noc2_valid;
wire tile_13_13_out_W_noc2_valid;
wire tile_13_13_out_N_noc2_yummy;
wire tile_13_13_out_S_noc2_yummy;
wire tile_13_13_out_E_noc2_yummy;
wire tile_13_13_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_13_13_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_13_13_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_13_13_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_13_13_out_W_noc3_data;
wire tile_13_13_out_N_noc3_valid;
wire tile_13_13_out_S_noc3_valid;
wire tile_13_13_out_E_noc3_valid;
wire tile_13_13_out_W_noc3_valid;
wire tile_13_13_out_N_noc3_yummy;
wire tile_13_13_out_S_noc3_yummy;
wire tile_13_13_out_E_noc3_yummy;
wire tile_13_13_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_14_13_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_14_13_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_14_13_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_14_13_out_W_noc1_data;
wire tile_14_13_out_N_noc1_valid;
wire tile_14_13_out_S_noc1_valid;
wire tile_14_13_out_E_noc1_valid;
wire tile_14_13_out_W_noc1_valid;
wire tile_14_13_out_N_noc1_yummy;
wire tile_14_13_out_S_noc1_yummy;
wire tile_14_13_out_E_noc1_yummy;
wire tile_14_13_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_14_13_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_14_13_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_14_13_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_14_13_out_W_noc2_data;
wire tile_14_13_out_N_noc2_valid;
wire tile_14_13_out_S_noc2_valid;
wire tile_14_13_out_E_noc2_valid;
wire tile_14_13_out_W_noc2_valid;
wire tile_14_13_out_N_noc2_yummy;
wire tile_14_13_out_S_noc2_yummy;
wire tile_14_13_out_E_noc2_yummy;
wire tile_14_13_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_14_13_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_14_13_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_14_13_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_14_13_out_W_noc3_data;
wire tile_14_13_out_N_noc3_valid;
wire tile_14_13_out_S_noc3_valid;
wire tile_14_13_out_E_noc3_valid;
wire tile_14_13_out_W_noc3_valid;
wire tile_14_13_out_N_noc3_yummy;
wire tile_14_13_out_S_noc3_yummy;
wire tile_14_13_out_E_noc3_yummy;
wire tile_14_13_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_15_13_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_15_13_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_15_13_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_15_13_out_W_noc1_data;
wire tile_15_13_out_N_noc1_valid;
wire tile_15_13_out_S_noc1_valid;
wire tile_15_13_out_E_noc1_valid;
wire tile_15_13_out_W_noc1_valid;
wire tile_15_13_out_N_noc1_yummy;
wire tile_15_13_out_S_noc1_yummy;
wire tile_15_13_out_E_noc1_yummy;
wire tile_15_13_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_15_13_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_15_13_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_15_13_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_15_13_out_W_noc2_data;
wire tile_15_13_out_N_noc2_valid;
wire tile_15_13_out_S_noc2_valid;
wire tile_15_13_out_E_noc2_valid;
wire tile_15_13_out_W_noc2_valid;
wire tile_15_13_out_N_noc2_yummy;
wire tile_15_13_out_S_noc2_yummy;
wire tile_15_13_out_E_noc2_yummy;
wire tile_15_13_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_15_13_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_15_13_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_15_13_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_15_13_out_W_noc3_data;
wire tile_15_13_out_N_noc3_valid;
wire tile_15_13_out_S_noc3_valid;
wire tile_15_13_out_E_noc3_valid;
wire tile_15_13_out_W_noc3_valid;
wire tile_15_13_out_N_noc3_yummy;
wire tile_15_13_out_S_noc3_yummy;
wire tile_15_13_out_E_noc3_yummy;
wire tile_15_13_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_0_14_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_0_14_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_0_14_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_0_14_out_W_noc1_data;
wire tile_0_14_out_N_noc1_valid;
wire tile_0_14_out_S_noc1_valid;
wire tile_0_14_out_E_noc1_valid;
wire tile_0_14_out_W_noc1_valid;
wire tile_0_14_out_N_noc1_yummy;
wire tile_0_14_out_S_noc1_yummy;
wire tile_0_14_out_E_noc1_yummy;
wire tile_0_14_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_0_14_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_0_14_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_0_14_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_0_14_out_W_noc2_data;
wire tile_0_14_out_N_noc2_valid;
wire tile_0_14_out_S_noc2_valid;
wire tile_0_14_out_E_noc2_valid;
wire tile_0_14_out_W_noc2_valid;
wire tile_0_14_out_N_noc2_yummy;
wire tile_0_14_out_S_noc2_yummy;
wire tile_0_14_out_E_noc2_yummy;
wire tile_0_14_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_0_14_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_0_14_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_0_14_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_0_14_out_W_noc3_data;
wire tile_0_14_out_N_noc3_valid;
wire tile_0_14_out_S_noc3_valid;
wire tile_0_14_out_E_noc3_valid;
wire tile_0_14_out_W_noc3_valid;
wire tile_0_14_out_N_noc3_yummy;
wire tile_0_14_out_S_noc3_yummy;
wire tile_0_14_out_E_noc3_yummy;
wire tile_0_14_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_1_14_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_1_14_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_1_14_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_1_14_out_W_noc1_data;
wire tile_1_14_out_N_noc1_valid;
wire tile_1_14_out_S_noc1_valid;
wire tile_1_14_out_E_noc1_valid;
wire tile_1_14_out_W_noc1_valid;
wire tile_1_14_out_N_noc1_yummy;
wire tile_1_14_out_S_noc1_yummy;
wire tile_1_14_out_E_noc1_yummy;
wire tile_1_14_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_1_14_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_1_14_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_1_14_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_1_14_out_W_noc2_data;
wire tile_1_14_out_N_noc2_valid;
wire tile_1_14_out_S_noc2_valid;
wire tile_1_14_out_E_noc2_valid;
wire tile_1_14_out_W_noc2_valid;
wire tile_1_14_out_N_noc2_yummy;
wire tile_1_14_out_S_noc2_yummy;
wire tile_1_14_out_E_noc2_yummy;
wire tile_1_14_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_1_14_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_1_14_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_1_14_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_1_14_out_W_noc3_data;
wire tile_1_14_out_N_noc3_valid;
wire tile_1_14_out_S_noc3_valid;
wire tile_1_14_out_E_noc3_valid;
wire tile_1_14_out_W_noc3_valid;
wire tile_1_14_out_N_noc3_yummy;
wire tile_1_14_out_S_noc3_yummy;
wire tile_1_14_out_E_noc3_yummy;
wire tile_1_14_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_2_14_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_2_14_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_2_14_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_2_14_out_W_noc1_data;
wire tile_2_14_out_N_noc1_valid;
wire tile_2_14_out_S_noc1_valid;
wire tile_2_14_out_E_noc1_valid;
wire tile_2_14_out_W_noc1_valid;
wire tile_2_14_out_N_noc1_yummy;
wire tile_2_14_out_S_noc1_yummy;
wire tile_2_14_out_E_noc1_yummy;
wire tile_2_14_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_2_14_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_2_14_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_2_14_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_2_14_out_W_noc2_data;
wire tile_2_14_out_N_noc2_valid;
wire tile_2_14_out_S_noc2_valid;
wire tile_2_14_out_E_noc2_valid;
wire tile_2_14_out_W_noc2_valid;
wire tile_2_14_out_N_noc2_yummy;
wire tile_2_14_out_S_noc2_yummy;
wire tile_2_14_out_E_noc2_yummy;
wire tile_2_14_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_2_14_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_2_14_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_2_14_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_2_14_out_W_noc3_data;
wire tile_2_14_out_N_noc3_valid;
wire tile_2_14_out_S_noc3_valid;
wire tile_2_14_out_E_noc3_valid;
wire tile_2_14_out_W_noc3_valid;
wire tile_2_14_out_N_noc3_yummy;
wire tile_2_14_out_S_noc3_yummy;
wire tile_2_14_out_E_noc3_yummy;
wire tile_2_14_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_3_14_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_3_14_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_3_14_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_3_14_out_W_noc1_data;
wire tile_3_14_out_N_noc1_valid;
wire tile_3_14_out_S_noc1_valid;
wire tile_3_14_out_E_noc1_valid;
wire tile_3_14_out_W_noc1_valid;
wire tile_3_14_out_N_noc1_yummy;
wire tile_3_14_out_S_noc1_yummy;
wire tile_3_14_out_E_noc1_yummy;
wire tile_3_14_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_3_14_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_3_14_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_3_14_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_3_14_out_W_noc2_data;
wire tile_3_14_out_N_noc2_valid;
wire tile_3_14_out_S_noc2_valid;
wire tile_3_14_out_E_noc2_valid;
wire tile_3_14_out_W_noc2_valid;
wire tile_3_14_out_N_noc2_yummy;
wire tile_3_14_out_S_noc2_yummy;
wire tile_3_14_out_E_noc2_yummy;
wire tile_3_14_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_3_14_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_3_14_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_3_14_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_3_14_out_W_noc3_data;
wire tile_3_14_out_N_noc3_valid;
wire tile_3_14_out_S_noc3_valid;
wire tile_3_14_out_E_noc3_valid;
wire tile_3_14_out_W_noc3_valid;
wire tile_3_14_out_N_noc3_yummy;
wire tile_3_14_out_S_noc3_yummy;
wire tile_3_14_out_E_noc3_yummy;
wire tile_3_14_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_4_14_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_4_14_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_4_14_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_4_14_out_W_noc1_data;
wire tile_4_14_out_N_noc1_valid;
wire tile_4_14_out_S_noc1_valid;
wire tile_4_14_out_E_noc1_valid;
wire tile_4_14_out_W_noc1_valid;
wire tile_4_14_out_N_noc1_yummy;
wire tile_4_14_out_S_noc1_yummy;
wire tile_4_14_out_E_noc1_yummy;
wire tile_4_14_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_4_14_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_4_14_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_4_14_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_4_14_out_W_noc2_data;
wire tile_4_14_out_N_noc2_valid;
wire tile_4_14_out_S_noc2_valid;
wire tile_4_14_out_E_noc2_valid;
wire tile_4_14_out_W_noc2_valid;
wire tile_4_14_out_N_noc2_yummy;
wire tile_4_14_out_S_noc2_yummy;
wire tile_4_14_out_E_noc2_yummy;
wire tile_4_14_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_4_14_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_4_14_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_4_14_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_4_14_out_W_noc3_data;
wire tile_4_14_out_N_noc3_valid;
wire tile_4_14_out_S_noc3_valid;
wire tile_4_14_out_E_noc3_valid;
wire tile_4_14_out_W_noc3_valid;
wire tile_4_14_out_N_noc3_yummy;
wire tile_4_14_out_S_noc3_yummy;
wire tile_4_14_out_E_noc3_yummy;
wire tile_4_14_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_5_14_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_5_14_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_5_14_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_5_14_out_W_noc1_data;
wire tile_5_14_out_N_noc1_valid;
wire tile_5_14_out_S_noc1_valid;
wire tile_5_14_out_E_noc1_valid;
wire tile_5_14_out_W_noc1_valid;
wire tile_5_14_out_N_noc1_yummy;
wire tile_5_14_out_S_noc1_yummy;
wire tile_5_14_out_E_noc1_yummy;
wire tile_5_14_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_5_14_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_5_14_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_5_14_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_5_14_out_W_noc2_data;
wire tile_5_14_out_N_noc2_valid;
wire tile_5_14_out_S_noc2_valid;
wire tile_5_14_out_E_noc2_valid;
wire tile_5_14_out_W_noc2_valid;
wire tile_5_14_out_N_noc2_yummy;
wire tile_5_14_out_S_noc2_yummy;
wire tile_5_14_out_E_noc2_yummy;
wire tile_5_14_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_5_14_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_5_14_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_5_14_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_5_14_out_W_noc3_data;
wire tile_5_14_out_N_noc3_valid;
wire tile_5_14_out_S_noc3_valid;
wire tile_5_14_out_E_noc3_valid;
wire tile_5_14_out_W_noc3_valid;
wire tile_5_14_out_N_noc3_yummy;
wire tile_5_14_out_S_noc3_yummy;
wire tile_5_14_out_E_noc3_yummy;
wire tile_5_14_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_6_14_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_6_14_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_6_14_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_6_14_out_W_noc1_data;
wire tile_6_14_out_N_noc1_valid;
wire tile_6_14_out_S_noc1_valid;
wire tile_6_14_out_E_noc1_valid;
wire tile_6_14_out_W_noc1_valid;
wire tile_6_14_out_N_noc1_yummy;
wire tile_6_14_out_S_noc1_yummy;
wire tile_6_14_out_E_noc1_yummy;
wire tile_6_14_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_6_14_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_6_14_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_6_14_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_6_14_out_W_noc2_data;
wire tile_6_14_out_N_noc2_valid;
wire tile_6_14_out_S_noc2_valid;
wire tile_6_14_out_E_noc2_valid;
wire tile_6_14_out_W_noc2_valid;
wire tile_6_14_out_N_noc2_yummy;
wire tile_6_14_out_S_noc2_yummy;
wire tile_6_14_out_E_noc2_yummy;
wire tile_6_14_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_6_14_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_6_14_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_6_14_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_6_14_out_W_noc3_data;
wire tile_6_14_out_N_noc3_valid;
wire tile_6_14_out_S_noc3_valid;
wire tile_6_14_out_E_noc3_valid;
wire tile_6_14_out_W_noc3_valid;
wire tile_6_14_out_N_noc3_yummy;
wire tile_6_14_out_S_noc3_yummy;
wire tile_6_14_out_E_noc3_yummy;
wire tile_6_14_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_7_14_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_7_14_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_7_14_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_7_14_out_W_noc1_data;
wire tile_7_14_out_N_noc1_valid;
wire tile_7_14_out_S_noc1_valid;
wire tile_7_14_out_E_noc1_valid;
wire tile_7_14_out_W_noc1_valid;
wire tile_7_14_out_N_noc1_yummy;
wire tile_7_14_out_S_noc1_yummy;
wire tile_7_14_out_E_noc1_yummy;
wire tile_7_14_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_7_14_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_7_14_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_7_14_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_7_14_out_W_noc2_data;
wire tile_7_14_out_N_noc2_valid;
wire tile_7_14_out_S_noc2_valid;
wire tile_7_14_out_E_noc2_valid;
wire tile_7_14_out_W_noc2_valid;
wire tile_7_14_out_N_noc2_yummy;
wire tile_7_14_out_S_noc2_yummy;
wire tile_7_14_out_E_noc2_yummy;
wire tile_7_14_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_7_14_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_7_14_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_7_14_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_7_14_out_W_noc3_data;
wire tile_7_14_out_N_noc3_valid;
wire tile_7_14_out_S_noc3_valid;
wire tile_7_14_out_E_noc3_valid;
wire tile_7_14_out_W_noc3_valid;
wire tile_7_14_out_N_noc3_yummy;
wire tile_7_14_out_S_noc3_yummy;
wire tile_7_14_out_E_noc3_yummy;
wire tile_7_14_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_8_14_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_8_14_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_8_14_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_8_14_out_W_noc1_data;
wire tile_8_14_out_N_noc1_valid;
wire tile_8_14_out_S_noc1_valid;
wire tile_8_14_out_E_noc1_valid;
wire tile_8_14_out_W_noc1_valid;
wire tile_8_14_out_N_noc1_yummy;
wire tile_8_14_out_S_noc1_yummy;
wire tile_8_14_out_E_noc1_yummy;
wire tile_8_14_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_8_14_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_8_14_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_8_14_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_8_14_out_W_noc2_data;
wire tile_8_14_out_N_noc2_valid;
wire tile_8_14_out_S_noc2_valid;
wire tile_8_14_out_E_noc2_valid;
wire tile_8_14_out_W_noc2_valid;
wire tile_8_14_out_N_noc2_yummy;
wire tile_8_14_out_S_noc2_yummy;
wire tile_8_14_out_E_noc2_yummy;
wire tile_8_14_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_8_14_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_8_14_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_8_14_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_8_14_out_W_noc3_data;
wire tile_8_14_out_N_noc3_valid;
wire tile_8_14_out_S_noc3_valid;
wire tile_8_14_out_E_noc3_valid;
wire tile_8_14_out_W_noc3_valid;
wire tile_8_14_out_N_noc3_yummy;
wire tile_8_14_out_S_noc3_yummy;
wire tile_8_14_out_E_noc3_yummy;
wire tile_8_14_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_9_14_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_9_14_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_9_14_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_9_14_out_W_noc1_data;
wire tile_9_14_out_N_noc1_valid;
wire tile_9_14_out_S_noc1_valid;
wire tile_9_14_out_E_noc1_valid;
wire tile_9_14_out_W_noc1_valid;
wire tile_9_14_out_N_noc1_yummy;
wire tile_9_14_out_S_noc1_yummy;
wire tile_9_14_out_E_noc1_yummy;
wire tile_9_14_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_9_14_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_9_14_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_9_14_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_9_14_out_W_noc2_data;
wire tile_9_14_out_N_noc2_valid;
wire tile_9_14_out_S_noc2_valid;
wire tile_9_14_out_E_noc2_valid;
wire tile_9_14_out_W_noc2_valid;
wire tile_9_14_out_N_noc2_yummy;
wire tile_9_14_out_S_noc2_yummy;
wire tile_9_14_out_E_noc2_yummy;
wire tile_9_14_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_9_14_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_9_14_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_9_14_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_9_14_out_W_noc3_data;
wire tile_9_14_out_N_noc3_valid;
wire tile_9_14_out_S_noc3_valid;
wire tile_9_14_out_E_noc3_valid;
wire tile_9_14_out_W_noc3_valid;
wire tile_9_14_out_N_noc3_yummy;
wire tile_9_14_out_S_noc3_yummy;
wire tile_9_14_out_E_noc3_yummy;
wire tile_9_14_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_10_14_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_10_14_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_10_14_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_10_14_out_W_noc1_data;
wire tile_10_14_out_N_noc1_valid;
wire tile_10_14_out_S_noc1_valid;
wire tile_10_14_out_E_noc1_valid;
wire tile_10_14_out_W_noc1_valid;
wire tile_10_14_out_N_noc1_yummy;
wire tile_10_14_out_S_noc1_yummy;
wire tile_10_14_out_E_noc1_yummy;
wire tile_10_14_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_10_14_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_10_14_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_10_14_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_10_14_out_W_noc2_data;
wire tile_10_14_out_N_noc2_valid;
wire tile_10_14_out_S_noc2_valid;
wire tile_10_14_out_E_noc2_valid;
wire tile_10_14_out_W_noc2_valid;
wire tile_10_14_out_N_noc2_yummy;
wire tile_10_14_out_S_noc2_yummy;
wire tile_10_14_out_E_noc2_yummy;
wire tile_10_14_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_10_14_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_10_14_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_10_14_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_10_14_out_W_noc3_data;
wire tile_10_14_out_N_noc3_valid;
wire tile_10_14_out_S_noc3_valid;
wire tile_10_14_out_E_noc3_valid;
wire tile_10_14_out_W_noc3_valid;
wire tile_10_14_out_N_noc3_yummy;
wire tile_10_14_out_S_noc3_yummy;
wire tile_10_14_out_E_noc3_yummy;
wire tile_10_14_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_11_14_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_11_14_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_11_14_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_11_14_out_W_noc1_data;
wire tile_11_14_out_N_noc1_valid;
wire tile_11_14_out_S_noc1_valid;
wire tile_11_14_out_E_noc1_valid;
wire tile_11_14_out_W_noc1_valid;
wire tile_11_14_out_N_noc1_yummy;
wire tile_11_14_out_S_noc1_yummy;
wire tile_11_14_out_E_noc1_yummy;
wire tile_11_14_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_11_14_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_11_14_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_11_14_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_11_14_out_W_noc2_data;
wire tile_11_14_out_N_noc2_valid;
wire tile_11_14_out_S_noc2_valid;
wire tile_11_14_out_E_noc2_valid;
wire tile_11_14_out_W_noc2_valid;
wire tile_11_14_out_N_noc2_yummy;
wire tile_11_14_out_S_noc2_yummy;
wire tile_11_14_out_E_noc2_yummy;
wire tile_11_14_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_11_14_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_11_14_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_11_14_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_11_14_out_W_noc3_data;
wire tile_11_14_out_N_noc3_valid;
wire tile_11_14_out_S_noc3_valid;
wire tile_11_14_out_E_noc3_valid;
wire tile_11_14_out_W_noc3_valid;
wire tile_11_14_out_N_noc3_yummy;
wire tile_11_14_out_S_noc3_yummy;
wire tile_11_14_out_E_noc3_yummy;
wire tile_11_14_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_12_14_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_12_14_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_12_14_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_12_14_out_W_noc1_data;
wire tile_12_14_out_N_noc1_valid;
wire tile_12_14_out_S_noc1_valid;
wire tile_12_14_out_E_noc1_valid;
wire tile_12_14_out_W_noc1_valid;
wire tile_12_14_out_N_noc1_yummy;
wire tile_12_14_out_S_noc1_yummy;
wire tile_12_14_out_E_noc1_yummy;
wire tile_12_14_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_12_14_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_12_14_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_12_14_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_12_14_out_W_noc2_data;
wire tile_12_14_out_N_noc2_valid;
wire tile_12_14_out_S_noc2_valid;
wire tile_12_14_out_E_noc2_valid;
wire tile_12_14_out_W_noc2_valid;
wire tile_12_14_out_N_noc2_yummy;
wire tile_12_14_out_S_noc2_yummy;
wire tile_12_14_out_E_noc2_yummy;
wire tile_12_14_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_12_14_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_12_14_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_12_14_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_12_14_out_W_noc3_data;
wire tile_12_14_out_N_noc3_valid;
wire tile_12_14_out_S_noc3_valid;
wire tile_12_14_out_E_noc3_valid;
wire tile_12_14_out_W_noc3_valid;
wire tile_12_14_out_N_noc3_yummy;
wire tile_12_14_out_S_noc3_yummy;
wire tile_12_14_out_E_noc3_yummy;
wire tile_12_14_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_13_14_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_13_14_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_13_14_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_13_14_out_W_noc1_data;
wire tile_13_14_out_N_noc1_valid;
wire tile_13_14_out_S_noc1_valid;
wire tile_13_14_out_E_noc1_valid;
wire tile_13_14_out_W_noc1_valid;
wire tile_13_14_out_N_noc1_yummy;
wire tile_13_14_out_S_noc1_yummy;
wire tile_13_14_out_E_noc1_yummy;
wire tile_13_14_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_13_14_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_13_14_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_13_14_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_13_14_out_W_noc2_data;
wire tile_13_14_out_N_noc2_valid;
wire tile_13_14_out_S_noc2_valid;
wire tile_13_14_out_E_noc2_valid;
wire tile_13_14_out_W_noc2_valid;
wire tile_13_14_out_N_noc2_yummy;
wire tile_13_14_out_S_noc2_yummy;
wire tile_13_14_out_E_noc2_yummy;
wire tile_13_14_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_13_14_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_13_14_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_13_14_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_13_14_out_W_noc3_data;
wire tile_13_14_out_N_noc3_valid;
wire tile_13_14_out_S_noc3_valid;
wire tile_13_14_out_E_noc3_valid;
wire tile_13_14_out_W_noc3_valid;
wire tile_13_14_out_N_noc3_yummy;
wire tile_13_14_out_S_noc3_yummy;
wire tile_13_14_out_E_noc3_yummy;
wire tile_13_14_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_14_14_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_14_14_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_14_14_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_14_14_out_W_noc1_data;
wire tile_14_14_out_N_noc1_valid;
wire tile_14_14_out_S_noc1_valid;
wire tile_14_14_out_E_noc1_valid;
wire tile_14_14_out_W_noc1_valid;
wire tile_14_14_out_N_noc1_yummy;
wire tile_14_14_out_S_noc1_yummy;
wire tile_14_14_out_E_noc1_yummy;
wire tile_14_14_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_14_14_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_14_14_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_14_14_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_14_14_out_W_noc2_data;
wire tile_14_14_out_N_noc2_valid;
wire tile_14_14_out_S_noc2_valid;
wire tile_14_14_out_E_noc2_valid;
wire tile_14_14_out_W_noc2_valid;
wire tile_14_14_out_N_noc2_yummy;
wire tile_14_14_out_S_noc2_yummy;
wire tile_14_14_out_E_noc2_yummy;
wire tile_14_14_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_14_14_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_14_14_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_14_14_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_14_14_out_W_noc3_data;
wire tile_14_14_out_N_noc3_valid;
wire tile_14_14_out_S_noc3_valid;
wire tile_14_14_out_E_noc3_valid;
wire tile_14_14_out_W_noc3_valid;
wire tile_14_14_out_N_noc3_yummy;
wire tile_14_14_out_S_noc3_yummy;
wire tile_14_14_out_E_noc3_yummy;
wire tile_14_14_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_15_14_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_15_14_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_15_14_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_15_14_out_W_noc1_data;
wire tile_15_14_out_N_noc1_valid;
wire tile_15_14_out_S_noc1_valid;
wire tile_15_14_out_E_noc1_valid;
wire tile_15_14_out_W_noc1_valid;
wire tile_15_14_out_N_noc1_yummy;
wire tile_15_14_out_S_noc1_yummy;
wire tile_15_14_out_E_noc1_yummy;
wire tile_15_14_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_15_14_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_15_14_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_15_14_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_15_14_out_W_noc2_data;
wire tile_15_14_out_N_noc2_valid;
wire tile_15_14_out_S_noc2_valid;
wire tile_15_14_out_E_noc2_valid;
wire tile_15_14_out_W_noc2_valid;
wire tile_15_14_out_N_noc2_yummy;
wire tile_15_14_out_S_noc2_yummy;
wire tile_15_14_out_E_noc2_yummy;
wire tile_15_14_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_15_14_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_15_14_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_15_14_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_15_14_out_W_noc3_data;
wire tile_15_14_out_N_noc3_valid;
wire tile_15_14_out_S_noc3_valid;
wire tile_15_14_out_E_noc3_valid;
wire tile_15_14_out_W_noc3_valid;
wire tile_15_14_out_N_noc3_yummy;
wire tile_15_14_out_S_noc3_yummy;
wire tile_15_14_out_E_noc3_yummy;
wire tile_15_14_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_0_15_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_0_15_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_0_15_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_0_15_out_W_noc1_data;
wire tile_0_15_out_N_noc1_valid;
wire tile_0_15_out_S_noc1_valid;
wire tile_0_15_out_E_noc1_valid;
wire tile_0_15_out_W_noc1_valid;
wire tile_0_15_out_N_noc1_yummy;
wire tile_0_15_out_S_noc1_yummy;
wire tile_0_15_out_E_noc1_yummy;
wire tile_0_15_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_0_15_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_0_15_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_0_15_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_0_15_out_W_noc2_data;
wire tile_0_15_out_N_noc2_valid;
wire tile_0_15_out_S_noc2_valid;
wire tile_0_15_out_E_noc2_valid;
wire tile_0_15_out_W_noc2_valid;
wire tile_0_15_out_N_noc2_yummy;
wire tile_0_15_out_S_noc2_yummy;
wire tile_0_15_out_E_noc2_yummy;
wire tile_0_15_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_0_15_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_0_15_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_0_15_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_0_15_out_W_noc3_data;
wire tile_0_15_out_N_noc3_valid;
wire tile_0_15_out_S_noc3_valid;
wire tile_0_15_out_E_noc3_valid;
wire tile_0_15_out_W_noc3_valid;
wire tile_0_15_out_N_noc3_yummy;
wire tile_0_15_out_S_noc3_yummy;
wire tile_0_15_out_E_noc3_yummy;
wire tile_0_15_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_1_15_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_1_15_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_1_15_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_1_15_out_W_noc1_data;
wire tile_1_15_out_N_noc1_valid;
wire tile_1_15_out_S_noc1_valid;
wire tile_1_15_out_E_noc1_valid;
wire tile_1_15_out_W_noc1_valid;
wire tile_1_15_out_N_noc1_yummy;
wire tile_1_15_out_S_noc1_yummy;
wire tile_1_15_out_E_noc1_yummy;
wire tile_1_15_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_1_15_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_1_15_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_1_15_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_1_15_out_W_noc2_data;
wire tile_1_15_out_N_noc2_valid;
wire tile_1_15_out_S_noc2_valid;
wire tile_1_15_out_E_noc2_valid;
wire tile_1_15_out_W_noc2_valid;
wire tile_1_15_out_N_noc2_yummy;
wire tile_1_15_out_S_noc2_yummy;
wire tile_1_15_out_E_noc2_yummy;
wire tile_1_15_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_1_15_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_1_15_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_1_15_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_1_15_out_W_noc3_data;
wire tile_1_15_out_N_noc3_valid;
wire tile_1_15_out_S_noc3_valid;
wire tile_1_15_out_E_noc3_valid;
wire tile_1_15_out_W_noc3_valid;
wire tile_1_15_out_N_noc3_yummy;
wire tile_1_15_out_S_noc3_yummy;
wire tile_1_15_out_E_noc3_yummy;
wire tile_1_15_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_2_15_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_2_15_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_2_15_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_2_15_out_W_noc1_data;
wire tile_2_15_out_N_noc1_valid;
wire tile_2_15_out_S_noc1_valid;
wire tile_2_15_out_E_noc1_valid;
wire tile_2_15_out_W_noc1_valid;
wire tile_2_15_out_N_noc1_yummy;
wire tile_2_15_out_S_noc1_yummy;
wire tile_2_15_out_E_noc1_yummy;
wire tile_2_15_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_2_15_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_2_15_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_2_15_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_2_15_out_W_noc2_data;
wire tile_2_15_out_N_noc2_valid;
wire tile_2_15_out_S_noc2_valid;
wire tile_2_15_out_E_noc2_valid;
wire tile_2_15_out_W_noc2_valid;
wire tile_2_15_out_N_noc2_yummy;
wire tile_2_15_out_S_noc2_yummy;
wire tile_2_15_out_E_noc2_yummy;
wire tile_2_15_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_2_15_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_2_15_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_2_15_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_2_15_out_W_noc3_data;
wire tile_2_15_out_N_noc3_valid;
wire tile_2_15_out_S_noc3_valid;
wire tile_2_15_out_E_noc3_valid;
wire tile_2_15_out_W_noc3_valid;
wire tile_2_15_out_N_noc3_yummy;
wire tile_2_15_out_S_noc3_yummy;
wire tile_2_15_out_E_noc3_yummy;
wire tile_2_15_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_3_15_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_3_15_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_3_15_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_3_15_out_W_noc1_data;
wire tile_3_15_out_N_noc1_valid;
wire tile_3_15_out_S_noc1_valid;
wire tile_3_15_out_E_noc1_valid;
wire tile_3_15_out_W_noc1_valid;
wire tile_3_15_out_N_noc1_yummy;
wire tile_3_15_out_S_noc1_yummy;
wire tile_3_15_out_E_noc1_yummy;
wire tile_3_15_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_3_15_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_3_15_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_3_15_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_3_15_out_W_noc2_data;
wire tile_3_15_out_N_noc2_valid;
wire tile_3_15_out_S_noc2_valid;
wire tile_3_15_out_E_noc2_valid;
wire tile_3_15_out_W_noc2_valid;
wire tile_3_15_out_N_noc2_yummy;
wire tile_3_15_out_S_noc2_yummy;
wire tile_3_15_out_E_noc2_yummy;
wire tile_3_15_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_3_15_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_3_15_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_3_15_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_3_15_out_W_noc3_data;
wire tile_3_15_out_N_noc3_valid;
wire tile_3_15_out_S_noc3_valid;
wire tile_3_15_out_E_noc3_valid;
wire tile_3_15_out_W_noc3_valid;
wire tile_3_15_out_N_noc3_yummy;
wire tile_3_15_out_S_noc3_yummy;
wire tile_3_15_out_E_noc3_yummy;
wire tile_3_15_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_4_15_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_4_15_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_4_15_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_4_15_out_W_noc1_data;
wire tile_4_15_out_N_noc1_valid;
wire tile_4_15_out_S_noc1_valid;
wire tile_4_15_out_E_noc1_valid;
wire tile_4_15_out_W_noc1_valid;
wire tile_4_15_out_N_noc1_yummy;
wire tile_4_15_out_S_noc1_yummy;
wire tile_4_15_out_E_noc1_yummy;
wire tile_4_15_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_4_15_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_4_15_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_4_15_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_4_15_out_W_noc2_data;
wire tile_4_15_out_N_noc2_valid;
wire tile_4_15_out_S_noc2_valid;
wire tile_4_15_out_E_noc2_valid;
wire tile_4_15_out_W_noc2_valid;
wire tile_4_15_out_N_noc2_yummy;
wire tile_4_15_out_S_noc2_yummy;
wire tile_4_15_out_E_noc2_yummy;
wire tile_4_15_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_4_15_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_4_15_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_4_15_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_4_15_out_W_noc3_data;
wire tile_4_15_out_N_noc3_valid;
wire tile_4_15_out_S_noc3_valid;
wire tile_4_15_out_E_noc3_valid;
wire tile_4_15_out_W_noc3_valid;
wire tile_4_15_out_N_noc3_yummy;
wire tile_4_15_out_S_noc3_yummy;
wire tile_4_15_out_E_noc3_yummy;
wire tile_4_15_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_5_15_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_5_15_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_5_15_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_5_15_out_W_noc1_data;
wire tile_5_15_out_N_noc1_valid;
wire tile_5_15_out_S_noc1_valid;
wire tile_5_15_out_E_noc1_valid;
wire tile_5_15_out_W_noc1_valid;
wire tile_5_15_out_N_noc1_yummy;
wire tile_5_15_out_S_noc1_yummy;
wire tile_5_15_out_E_noc1_yummy;
wire tile_5_15_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_5_15_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_5_15_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_5_15_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_5_15_out_W_noc2_data;
wire tile_5_15_out_N_noc2_valid;
wire tile_5_15_out_S_noc2_valid;
wire tile_5_15_out_E_noc2_valid;
wire tile_5_15_out_W_noc2_valid;
wire tile_5_15_out_N_noc2_yummy;
wire tile_5_15_out_S_noc2_yummy;
wire tile_5_15_out_E_noc2_yummy;
wire tile_5_15_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_5_15_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_5_15_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_5_15_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_5_15_out_W_noc3_data;
wire tile_5_15_out_N_noc3_valid;
wire tile_5_15_out_S_noc3_valid;
wire tile_5_15_out_E_noc3_valid;
wire tile_5_15_out_W_noc3_valid;
wire tile_5_15_out_N_noc3_yummy;
wire tile_5_15_out_S_noc3_yummy;
wire tile_5_15_out_E_noc3_yummy;
wire tile_5_15_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_6_15_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_6_15_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_6_15_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_6_15_out_W_noc1_data;
wire tile_6_15_out_N_noc1_valid;
wire tile_6_15_out_S_noc1_valid;
wire tile_6_15_out_E_noc1_valid;
wire tile_6_15_out_W_noc1_valid;
wire tile_6_15_out_N_noc1_yummy;
wire tile_6_15_out_S_noc1_yummy;
wire tile_6_15_out_E_noc1_yummy;
wire tile_6_15_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_6_15_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_6_15_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_6_15_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_6_15_out_W_noc2_data;
wire tile_6_15_out_N_noc2_valid;
wire tile_6_15_out_S_noc2_valid;
wire tile_6_15_out_E_noc2_valid;
wire tile_6_15_out_W_noc2_valid;
wire tile_6_15_out_N_noc2_yummy;
wire tile_6_15_out_S_noc2_yummy;
wire tile_6_15_out_E_noc2_yummy;
wire tile_6_15_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_6_15_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_6_15_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_6_15_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_6_15_out_W_noc3_data;
wire tile_6_15_out_N_noc3_valid;
wire tile_6_15_out_S_noc3_valid;
wire tile_6_15_out_E_noc3_valid;
wire tile_6_15_out_W_noc3_valid;
wire tile_6_15_out_N_noc3_yummy;
wire tile_6_15_out_S_noc3_yummy;
wire tile_6_15_out_E_noc3_yummy;
wire tile_6_15_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_7_15_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_7_15_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_7_15_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_7_15_out_W_noc1_data;
wire tile_7_15_out_N_noc1_valid;
wire tile_7_15_out_S_noc1_valid;
wire tile_7_15_out_E_noc1_valid;
wire tile_7_15_out_W_noc1_valid;
wire tile_7_15_out_N_noc1_yummy;
wire tile_7_15_out_S_noc1_yummy;
wire tile_7_15_out_E_noc1_yummy;
wire tile_7_15_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_7_15_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_7_15_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_7_15_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_7_15_out_W_noc2_data;
wire tile_7_15_out_N_noc2_valid;
wire tile_7_15_out_S_noc2_valid;
wire tile_7_15_out_E_noc2_valid;
wire tile_7_15_out_W_noc2_valid;
wire tile_7_15_out_N_noc2_yummy;
wire tile_7_15_out_S_noc2_yummy;
wire tile_7_15_out_E_noc2_yummy;
wire tile_7_15_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_7_15_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_7_15_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_7_15_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_7_15_out_W_noc3_data;
wire tile_7_15_out_N_noc3_valid;
wire tile_7_15_out_S_noc3_valid;
wire tile_7_15_out_E_noc3_valid;
wire tile_7_15_out_W_noc3_valid;
wire tile_7_15_out_N_noc3_yummy;
wire tile_7_15_out_S_noc3_yummy;
wire tile_7_15_out_E_noc3_yummy;
wire tile_7_15_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_8_15_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_8_15_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_8_15_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_8_15_out_W_noc1_data;
wire tile_8_15_out_N_noc1_valid;
wire tile_8_15_out_S_noc1_valid;
wire tile_8_15_out_E_noc1_valid;
wire tile_8_15_out_W_noc1_valid;
wire tile_8_15_out_N_noc1_yummy;
wire tile_8_15_out_S_noc1_yummy;
wire tile_8_15_out_E_noc1_yummy;
wire tile_8_15_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_8_15_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_8_15_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_8_15_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_8_15_out_W_noc2_data;
wire tile_8_15_out_N_noc2_valid;
wire tile_8_15_out_S_noc2_valid;
wire tile_8_15_out_E_noc2_valid;
wire tile_8_15_out_W_noc2_valid;
wire tile_8_15_out_N_noc2_yummy;
wire tile_8_15_out_S_noc2_yummy;
wire tile_8_15_out_E_noc2_yummy;
wire tile_8_15_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_8_15_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_8_15_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_8_15_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_8_15_out_W_noc3_data;
wire tile_8_15_out_N_noc3_valid;
wire tile_8_15_out_S_noc3_valid;
wire tile_8_15_out_E_noc3_valid;
wire tile_8_15_out_W_noc3_valid;
wire tile_8_15_out_N_noc3_yummy;
wire tile_8_15_out_S_noc3_yummy;
wire tile_8_15_out_E_noc3_yummy;
wire tile_8_15_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_9_15_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_9_15_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_9_15_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_9_15_out_W_noc1_data;
wire tile_9_15_out_N_noc1_valid;
wire tile_9_15_out_S_noc1_valid;
wire tile_9_15_out_E_noc1_valid;
wire tile_9_15_out_W_noc1_valid;
wire tile_9_15_out_N_noc1_yummy;
wire tile_9_15_out_S_noc1_yummy;
wire tile_9_15_out_E_noc1_yummy;
wire tile_9_15_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_9_15_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_9_15_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_9_15_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_9_15_out_W_noc2_data;
wire tile_9_15_out_N_noc2_valid;
wire tile_9_15_out_S_noc2_valid;
wire tile_9_15_out_E_noc2_valid;
wire tile_9_15_out_W_noc2_valid;
wire tile_9_15_out_N_noc2_yummy;
wire tile_9_15_out_S_noc2_yummy;
wire tile_9_15_out_E_noc2_yummy;
wire tile_9_15_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_9_15_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_9_15_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_9_15_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_9_15_out_W_noc3_data;
wire tile_9_15_out_N_noc3_valid;
wire tile_9_15_out_S_noc3_valid;
wire tile_9_15_out_E_noc3_valid;
wire tile_9_15_out_W_noc3_valid;
wire tile_9_15_out_N_noc3_yummy;
wire tile_9_15_out_S_noc3_yummy;
wire tile_9_15_out_E_noc3_yummy;
wire tile_9_15_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_10_15_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_10_15_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_10_15_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_10_15_out_W_noc1_data;
wire tile_10_15_out_N_noc1_valid;
wire tile_10_15_out_S_noc1_valid;
wire tile_10_15_out_E_noc1_valid;
wire tile_10_15_out_W_noc1_valid;
wire tile_10_15_out_N_noc1_yummy;
wire tile_10_15_out_S_noc1_yummy;
wire tile_10_15_out_E_noc1_yummy;
wire tile_10_15_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_10_15_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_10_15_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_10_15_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_10_15_out_W_noc2_data;
wire tile_10_15_out_N_noc2_valid;
wire tile_10_15_out_S_noc2_valid;
wire tile_10_15_out_E_noc2_valid;
wire tile_10_15_out_W_noc2_valid;
wire tile_10_15_out_N_noc2_yummy;
wire tile_10_15_out_S_noc2_yummy;
wire tile_10_15_out_E_noc2_yummy;
wire tile_10_15_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_10_15_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_10_15_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_10_15_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_10_15_out_W_noc3_data;
wire tile_10_15_out_N_noc3_valid;
wire tile_10_15_out_S_noc3_valid;
wire tile_10_15_out_E_noc3_valid;
wire tile_10_15_out_W_noc3_valid;
wire tile_10_15_out_N_noc3_yummy;
wire tile_10_15_out_S_noc3_yummy;
wire tile_10_15_out_E_noc3_yummy;
wire tile_10_15_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_11_15_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_11_15_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_11_15_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_11_15_out_W_noc1_data;
wire tile_11_15_out_N_noc1_valid;
wire tile_11_15_out_S_noc1_valid;
wire tile_11_15_out_E_noc1_valid;
wire tile_11_15_out_W_noc1_valid;
wire tile_11_15_out_N_noc1_yummy;
wire tile_11_15_out_S_noc1_yummy;
wire tile_11_15_out_E_noc1_yummy;
wire tile_11_15_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_11_15_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_11_15_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_11_15_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_11_15_out_W_noc2_data;
wire tile_11_15_out_N_noc2_valid;
wire tile_11_15_out_S_noc2_valid;
wire tile_11_15_out_E_noc2_valid;
wire tile_11_15_out_W_noc2_valid;
wire tile_11_15_out_N_noc2_yummy;
wire tile_11_15_out_S_noc2_yummy;
wire tile_11_15_out_E_noc2_yummy;
wire tile_11_15_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_11_15_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_11_15_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_11_15_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_11_15_out_W_noc3_data;
wire tile_11_15_out_N_noc3_valid;
wire tile_11_15_out_S_noc3_valid;
wire tile_11_15_out_E_noc3_valid;
wire tile_11_15_out_W_noc3_valid;
wire tile_11_15_out_N_noc3_yummy;
wire tile_11_15_out_S_noc3_yummy;
wire tile_11_15_out_E_noc3_yummy;
wire tile_11_15_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_12_15_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_12_15_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_12_15_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_12_15_out_W_noc1_data;
wire tile_12_15_out_N_noc1_valid;
wire tile_12_15_out_S_noc1_valid;
wire tile_12_15_out_E_noc1_valid;
wire tile_12_15_out_W_noc1_valid;
wire tile_12_15_out_N_noc1_yummy;
wire tile_12_15_out_S_noc1_yummy;
wire tile_12_15_out_E_noc1_yummy;
wire tile_12_15_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_12_15_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_12_15_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_12_15_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_12_15_out_W_noc2_data;
wire tile_12_15_out_N_noc2_valid;
wire tile_12_15_out_S_noc2_valid;
wire tile_12_15_out_E_noc2_valid;
wire tile_12_15_out_W_noc2_valid;
wire tile_12_15_out_N_noc2_yummy;
wire tile_12_15_out_S_noc2_yummy;
wire tile_12_15_out_E_noc2_yummy;
wire tile_12_15_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_12_15_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_12_15_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_12_15_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_12_15_out_W_noc3_data;
wire tile_12_15_out_N_noc3_valid;
wire tile_12_15_out_S_noc3_valid;
wire tile_12_15_out_E_noc3_valid;
wire tile_12_15_out_W_noc3_valid;
wire tile_12_15_out_N_noc3_yummy;
wire tile_12_15_out_S_noc3_yummy;
wire tile_12_15_out_E_noc3_yummy;
wire tile_12_15_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_13_15_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_13_15_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_13_15_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_13_15_out_W_noc1_data;
wire tile_13_15_out_N_noc1_valid;
wire tile_13_15_out_S_noc1_valid;
wire tile_13_15_out_E_noc1_valid;
wire tile_13_15_out_W_noc1_valid;
wire tile_13_15_out_N_noc1_yummy;
wire tile_13_15_out_S_noc1_yummy;
wire tile_13_15_out_E_noc1_yummy;
wire tile_13_15_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_13_15_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_13_15_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_13_15_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_13_15_out_W_noc2_data;
wire tile_13_15_out_N_noc2_valid;
wire tile_13_15_out_S_noc2_valid;
wire tile_13_15_out_E_noc2_valid;
wire tile_13_15_out_W_noc2_valid;
wire tile_13_15_out_N_noc2_yummy;
wire tile_13_15_out_S_noc2_yummy;
wire tile_13_15_out_E_noc2_yummy;
wire tile_13_15_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_13_15_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_13_15_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_13_15_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_13_15_out_W_noc3_data;
wire tile_13_15_out_N_noc3_valid;
wire tile_13_15_out_S_noc3_valid;
wire tile_13_15_out_E_noc3_valid;
wire tile_13_15_out_W_noc3_valid;
wire tile_13_15_out_N_noc3_yummy;
wire tile_13_15_out_S_noc3_yummy;
wire tile_13_15_out_E_noc3_yummy;
wire tile_13_15_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_14_15_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_14_15_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_14_15_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_14_15_out_W_noc1_data;
wire tile_14_15_out_N_noc1_valid;
wire tile_14_15_out_S_noc1_valid;
wire tile_14_15_out_E_noc1_valid;
wire tile_14_15_out_W_noc1_valid;
wire tile_14_15_out_N_noc1_yummy;
wire tile_14_15_out_S_noc1_yummy;
wire tile_14_15_out_E_noc1_yummy;
wire tile_14_15_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_14_15_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_14_15_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_14_15_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_14_15_out_W_noc2_data;
wire tile_14_15_out_N_noc2_valid;
wire tile_14_15_out_S_noc2_valid;
wire tile_14_15_out_E_noc2_valid;
wire tile_14_15_out_W_noc2_valid;
wire tile_14_15_out_N_noc2_yummy;
wire tile_14_15_out_S_noc2_yummy;
wire tile_14_15_out_E_noc2_yummy;
wire tile_14_15_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_14_15_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_14_15_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_14_15_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_14_15_out_W_noc3_data;
wire tile_14_15_out_N_noc3_valid;
wire tile_14_15_out_S_noc3_valid;
wire tile_14_15_out_E_noc3_valid;
wire tile_14_15_out_W_noc3_valid;
wire tile_14_15_out_N_noc3_yummy;
wire tile_14_15_out_S_noc3_yummy;
wire tile_14_15_out_E_noc3_yummy;
wire tile_14_15_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] tile_15_15_out_N_noc1_data;
wire [`DATA_WIDTH-1:0] tile_15_15_out_S_noc1_data;
wire [`DATA_WIDTH-1:0] tile_15_15_out_E_noc1_data;
wire [`DATA_WIDTH-1:0] tile_15_15_out_W_noc1_data;
wire tile_15_15_out_N_noc1_valid;
wire tile_15_15_out_S_noc1_valid;
wire tile_15_15_out_E_noc1_valid;
wire tile_15_15_out_W_noc1_valid;
wire tile_15_15_out_N_noc1_yummy;
wire tile_15_15_out_S_noc1_yummy;
wire tile_15_15_out_E_noc1_yummy;
wire tile_15_15_out_W_noc1_yummy;
wire [`DATA_WIDTH-1:0] tile_15_15_out_N_noc2_data;
wire [`DATA_WIDTH-1:0] tile_15_15_out_S_noc2_data;
wire [`DATA_WIDTH-1:0] tile_15_15_out_E_noc2_data;
wire [`DATA_WIDTH-1:0] tile_15_15_out_W_noc2_data;
wire tile_15_15_out_N_noc2_valid;
wire tile_15_15_out_S_noc2_valid;
wire tile_15_15_out_E_noc2_valid;
wire tile_15_15_out_W_noc2_valid;
wire tile_15_15_out_N_noc2_yummy;
wire tile_15_15_out_S_noc2_yummy;
wire tile_15_15_out_E_noc2_yummy;
wire tile_15_15_out_W_noc2_yummy;
wire [`DATA_WIDTH-1:0] tile_15_15_out_N_noc3_data;
wire [`DATA_WIDTH-1:0] tile_15_15_out_S_noc3_data;
wire [`DATA_WIDTH-1:0] tile_15_15_out_E_noc3_data;
wire [`DATA_WIDTH-1:0] tile_15_15_out_W_noc3_data;
wire tile_15_15_out_N_noc3_valid;
wire tile_15_15_out_S_noc3_valid;
wire tile_15_15_out_E_noc3_valid;
wire tile_15_15_out_W_noc3_valid;
wire tile_15_15_out_N_noc3_yummy;
wire tile_15_15_out_S_noc3_yummy;
wire tile_15_15_out_E_noc3_yummy;
wire tile_15_15_out_W_noc3_yummy;
wire [`DATA_WIDTH-1:0] dummy_out_N_noc1_data = `DATA_WIDTH'b0;
wire [`DATA_WIDTH-1:0] dummy_out_S_noc1_data = `DATA_WIDTH'b0;
wire [`DATA_WIDTH-1:0] dummy_out_E_noc1_data = `DATA_WIDTH'b0;
wire [`DATA_WIDTH-1:0] dummy_out_W_noc1_data = `DATA_WIDTH'b0;
wire dummy_out_N_noc1_valid = 1'b0;
wire dummy_out_S_noc1_valid = 1'b0;
wire dummy_out_E_noc1_valid = 1'b0;
wire dummy_out_W_noc1_valid = 1'b0;
wire dummy_out_N_noc1_yummy = 1'b0;
wire dummy_out_S_noc1_yummy = 1'b0;
wire dummy_out_E_noc1_yummy = 1'b0;
wire dummy_out_W_noc1_yummy = 1'b0;
wire [`DATA_WIDTH-1:0] dummy_out_N_noc2_data = `DATA_WIDTH'b0;
wire [`DATA_WIDTH-1:0] dummy_out_S_noc2_data = `DATA_WIDTH'b0;
wire [`DATA_WIDTH-1:0] dummy_out_E_noc2_data = `DATA_WIDTH'b0;
wire [`DATA_WIDTH-1:0] dummy_out_W_noc2_data = `DATA_WIDTH'b0;
wire dummy_out_N_noc2_valid = 1'b0;
wire dummy_out_S_noc2_valid = 1'b0;
wire dummy_out_E_noc2_valid = 1'b0;
wire dummy_out_W_noc2_valid = 1'b0;
wire dummy_out_N_noc2_yummy = 1'b0;
wire dummy_out_S_noc2_yummy = 1'b0;
wire dummy_out_E_noc2_yummy = 1'b0;
wire dummy_out_W_noc2_yummy = 1'b0;
wire [`DATA_WIDTH-1:0] dummy_out_N_noc3_data = `DATA_WIDTH'b0;
wire [`DATA_WIDTH-1:0] dummy_out_S_noc3_data = `DATA_WIDTH'b0;
wire [`DATA_WIDTH-1:0] dummy_out_E_noc3_data = `DATA_WIDTH'b0;
wire [`DATA_WIDTH-1:0] dummy_out_W_noc3_data = `DATA_WIDTH'b0;
wire dummy_out_N_noc3_valid = 1'b0;
wire dummy_out_S_noc3_valid = 1'b0;
wire dummy_out_E_noc3_valid = 1'b0;
wire dummy_out_W_noc3_valid = 1'b0;
wire dummy_out_N_noc3_yummy = 1'b0;
wire dummy_out_S_noc3_yummy = 1'b0;
wire dummy_out_E_noc3_yummy = 1'b0;
wire dummy_out_W_noc3_yummy = 1'b0;
wire [`DATA_WIDTH-1:0] offchip_out_E_noc1_data;
wire offchip_out_E_noc1_valid;
wire offchip_out_E_noc1_yummy;
wire [`DATA_WIDTH-1:0] offchip_out_E_noc2_data;
wire offchip_out_E_noc2_valid;
wire offchip_out_E_noc2_yummy;
wire [`DATA_WIDTH-1:0] offchip_out_E_noc3_data;
wire offchip_out_E_noc3_valid;
wire offchip_out_E_noc3_yummy;


   //////////////////////
   // Sequential logic
   //////////////////////

   // trin 2/3/15:
   // rst in the tile is flopped for an additional cycle
   // we'll do the same for all other modules at the chip.v level
   always @ (posedge clk_muxed)
      rst_n_inter_sync_f <= rst_n_inter_sync;

   always @ (posedge io_clk_inter)
      io_clk_rst_n_inter_sync_f <= io_clk_rst_n_inter_sync;

`ifndef PITON_NO_CHIP_BRIDGE
   // Buffer chip bridge inputs
   always @(posedge io_clk_inter)
   begin
`ifdef PITON_PROTO
       if(~io_clk_rst_n_inter_sync_f)
`else // ifndef PITON_PROTO
       if(~rst_n_inter_sync_f)
`endif
       begin
           intf_chip_data_inter_buf_f <= 0;
           intf_chip_channel_inter_buf_f <= 0;
           chip_intf_credit_back_inter_buf_f <= 0;
       end
       else
       begin
           intf_chip_data_inter_buf_f <= intf_chip_data_inter;
           intf_chip_channel_inter_buf_f <= intf_chip_channel_inter;
           chip_intf_credit_back_inter_buf_f <= chip_intf_credit_back_inter;
       end
   end
`endif // endif PITON_NO_CHIP_BRIDGE

   ////////////////////////
   // Combinational Logic
   ////////////////////////

   // Need to assign missing inputs and outputs if synthesizing
   // chip for FPGA standalone
`ifdef PITON_CHIP_FPGA
   assign slew = 1'b1;
   assign impsel1 = 1'b1;
   assign impsel2 = 1'b1;

   assign pll_rst_n = 1'b1;

   assign clk_en = 1'b1;

   assign pll_lock = 1'b1;
   assign pll_bypass = 1'b1;
   assign pll_rangea = 5'b0;

   assign clk_mux_sel = 2'b0;

   assign jtag_clk = 1'b0;
   assign jtag_rst_l = 1'b1;
   assign jtag_modesel = 1'b1;
   assign jtag_datain = 1'b0;

   assign async_mux = 1'b1;

   assign oram_on = 1'b0;
   assign oram_traffic_gen = 1'b0;
   assign oram_dummy_gen = 1'b0;

   assign piton_prsnt_n = ~rst_n_inter_sync;
   assign piton_ready_n = ~rst_n_inter_sync;

`ifdef PITON_FPGA_CLKS_GEN
   assign leds[0] = mmcm_locked;
`else // ifndef PITON_FPGA_CLKS_GEN
   assign leds[0] = 1'b1;
`endif // endif PITON_FPGA_CLKS_GEN
   assign leds[1] = rst_n_inter_sync;
   assign leds[2] = io_clk_rst_n_inter_sync;
   assign leds[3] = processor_offchip_noc1_valid;
   assign leds[4] = processor_offchip_noc2_valid;
   assign leds[5] = offchip_processor_noc2_valid;
   assign leds[6] = offchip_processor_noc3_valid;
   assign leds[7] = 1'b0;

`endif // endif PITON_CHIP_FPGA

   // Connecting chip_bridge data to tiles/ORAM

assign proc_oram_valid = tile_0_0_out_W_noc2_valid;
assign proc_oram_data = tile_0_0_out_W_noc2_data;
assign oram_proc_yummy = tile_0_0_out_W_noc3_yummy;

   assign offchip_oram_valid = offchip_processor_noc3_valid;
   assign offchip_oram_data = offchip_processor_noc3_data;
   assign oram_offchip_yummy = processor_offchip_noc2_yummy;

assign processor_offchip_noc1_valid = tile_0_0_out_W_noc1_valid;
assign processor_offchip_noc1_data = tile_0_0_out_W_noc1_data;
assign offchip_processor_noc1_yummy = tile_0_0_out_W_noc1_yummy;

   assign processor_offchip_noc2_valid = oram_offchip_valid;
   assign processor_offchip_noc2_data = oram_offchip_data;

assign offchip_processor_noc2_yummy = tile_0_0_out_W_noc2_yummy;
assign processor_offchip_noc3_valid = tile_0_0_out_W_noc3_valid;
assign processor_offchip_noc3_data = tile_0_0_out_W_noc3_data;

   assign offchip_processor_noc3_yummy = offchip_oram_yummy;

assign offchip_out_E_noc1_data = offchip_processor_noc1_data;
assign offchip_out_E_noc1_valid = offchip_processor_noc1_valid;
assign offchip_out_E_noc1_yummy = processor_offchip_noc1_yummy;
assign offchip_out_E_noc2_data = offchip_processor_noc2_data;
assign offchip_out_E_noc2_valid = offchip_processor_noc2_valid;
assign offchip_out_E_noc2_yummy = proc_oram_yummy; //going to processor
assign offchip_out_E_noc3_data = oram_proc_data;
assign offchip_out_E_noc3_valid = oram_proc_valid;
assign offchip_out_E_noc3_yummy = processor_offchip_noc3_yummy;


   // trin: off-chip channel mux when disabling oram
   always @ *
   begin
     // default is bypassing
     oram_offchip_valid = proc_oram_valid;
     oram_offchip_data = proc_oram_data;
     proc_oram_yummy = oram_offchip_yummy;
     oram_proc_valid = offchip_oram_valid;
     oram_proc_data = offchip_oram_data;
     offchip_oram_yummy = oram_proc_yummy;

     if (oram_on_inter)
     begin
       oram_offchip_valid = oram_offchip_valid_oram;
       oram_offchip_data = oram_offchip_data_oram;
       proc_oram_yummy = proc_oram_yummy_oram;
       oram_proc_valid = oram_proc_valid_oram;
       oram_proc_data = oram_proc_data_oram;
       offchip_oram_yummy = offchip_oram_yummy_oram;
     end
   end

   // Merge all JTAG outputs from tiles together
assign tiles_jtag_ucb_val = tile0_jtag_ucb_val | tile16_jtag_ucb_val | tile32_jtag_ucb_val | tile48_jtag_ucb_val | tile64_jtag_ucb_val | tile80_jtag_ucb_val | tile96_jtag_ucb_val | tile112_jtag_ucb_val | tile128_jtag_ucb_val | tile144_jtag_ucb_val | tile160_jtag_ucb_val | tile176_jtag_ucb_val | tile192_jtag_ucb_val | tile208_jtag_ucb_val | tile224_jtag_ucb_val | tile240_jtag_ucb_val | tile1_jtag_ucb_val | tile17_jtag_ucb_val | tile33_jtag_ucb_val | tile49_jtag_ucb_val | tile65_jtag_ucb_val | tile81_jtag_ucb_val | tile97_jtag_ucb_val | tile113_jtag_ucb_val | tile129_jtag_ucb_val | tile145_jtag_ucb_val | tile161_jtag_ucb_val | tile177_jtag_ucb_val | tile193_jtag_ucb_val | tile209_jtag_ucb_val | tile225_jtag_ucb_val | tile241_jtag_ucb_val | tile2_jtag_ucb_val | tile18_jtag_ucb_val | tile34_jtag_ucb_val | tile50_jtag_ucb_val | tile66_jtag_ucb_val | tile82_jtag_ucb_val | tile98_jtag_ucb_val | tile114_jtag_ucb_val | tile130_jtag_ucb_val | tile146_jtag_ucb_val | tile162_jtag_ucb_val | tile178_jtag_ucb_val | tile194_jtag_ucb_val | tile210_jtag_ucb_val | tile226_jtag_ucb_val | tile242_jtag_ucb_val | tile3_jtag_ucb_val | tile19_jtag_ucb_val | tile35_jtag_ucb_val | tile51_jtag_ucb_val | tile67_jtag_ucb_val | tile83_jtag_ucb_val | tile99_jtag_ucb_val | tile115_jtag_ucb_val | tile131_jtag_ucb_val | tile147_jtag_ucb_val | tile163_jtag_ucb_val | tile179_jtag_ucb_val | tile195_jtag_ucb_val | tile211_jtag_ucb_val | tile227_jtag_ucb_val | tile243_jtag_ucb_val | tile4_jtag_ucb_val | tile20_jtag_ucb_val | tile36_jtag_ucb_val | tile52_jtag_ucb_val | tile68_jtag_ucb_val | tile84_jtag_ucb_val | tile100_jtag_ucb_val | tile116_jtag_ucb_val | tile132_jtag_ucb_val | tile148_jtag_ucb_val | tile164_jtag_ucb_val | tile180_jtag_ucb_val | tile196_jtag_ucb_val | tile212_jtag_ucb_val | tile228_jtag_ucb_val | tile244_jtag_ucb_val | tile5_jtag_ucb_val | tile21_jtag_ucb_val | tile37_jtag_ucb_val | tile53_jtag_ucb_val | tile69_jtag_ucb_val | tile85_jtag_ucb_val | tile101_jtag_ucb_val | tile117_jtag_ucb_val | tile133_jtag_ucb_val | tile149_jtag_ucb_val | tile165_jtag_ucb_val | tile181_jtag_ucb_val | tile197_jtag_ucb_val | tile213_jtag_ucb_val | tile229_jtag_ucb_val | tile245_jtag_ucb_val | tile6_jtag_ucb_val | tile22_jtag_ucb_val | tile38_jtag_ucb_val | tile54_jtag_ucb_val | tile70_jtag_ucb_val | tile86_jtag_ucb_val | tile102_jtag_ucb_val | tile118_jtag_ucb_val | tile134_jtag_ucb_val | tile150_jtag_ucb_val | tile166_jtag_ucb_val | tile182_jtag_ucb_val | tile198_jtag_ucb_val | tile214_jtag_ucb_val | tile230_jtag_ucb_val | tile246_jtag_ucb_val | tile7_jtag_ucb_val | tile23_jtag_ucb_val | tile39_jtag_ucb_val | tile55_jtag_ucb_val | tile71_jtag_ucb_val | tile87_jtag_ucb_val | tile103_jtag_ucb_val | tile119_jtag_ucb_val | tile135_jtag_ucb_val | tile151_jtag_ucb_val | tile167_jtag_ucb_val | tile183_jtag_ucb_val | tile199_jtag_ucb_val | tile215_jtag_ucb_val | tile231_jtag_ucb_val | tile247_jtag_ucb_val | tile8_jtag_ucb_val | tile24_jtag_ucb_val | tile40_jtag_ucb_val | tile56_jtag_ucb_val | tile72_jtag_ucb_val | tile88_jtag_ucb_val | tile104_jtag_ucb_val | tile120_jtag_ucb_val | tile136_jtag_ucb_val | tile152_jtag_ucb_val | tile168_jtag_ucb_val | tile184_jtag_ucb_val | tile200_jtag_ucb_val | tile216_jtag_ucb_val | tile232_jtag_ucb_val | tile248_jtag_ucb_val | tile9_jtag_ucb_val | tile25_jtag_ucb_val | tile41_jtag_ucb_val | tile57_jtag_ucb_val | tile73_jtag_ucb_val | tile89_jtag_ucb_val | tile105_jtag_ucb_val | tile121_jtag_ucb_val | tile137_jtag_ucb_val | tile153_jtag_ucb_val | tile169_jtag_ucb_val | tile185_jtag_ucb_val | tile201_jtag_ucb_val | tile217_jtag_ucb_val | tile233_jtag_ucb_val | tile249_jtag_ucb_val | tile10_jtag_ucb_val | tile26_jtag_ucb_val | tile42_jtag_ucb_val | tile58_jtag_ucb_val | tile74_jtag_ucb_val | tile90_jtag_ucb_val | tile106_jtag_ucb_val | tile122_jtag_ucb_val | tile138_jtag_ucb_val | tile154_jtag_ucb_val | tile170_jtag_ucb_val | tile186_jtag_ucb_val | tile202_jtag_ucb_val | tile218_jtag_ucb_val | tile234_jtag_ucb_val | tile250_jtag_ucb_val | tile11_jtag_ucb_val | tile27_jtag_ucb_val | tile43_jtag_ucb_val | tile59_jtag_ucb_val | tile75_jtag_ucb_val | tile91_jtag_ucb_val | tile107_jtag_ucb_val | tile123_jtag_ucb_val | tile139_jtag_ucb_val | tile155_jtag_ucb_val | tile171_jtag_ucb_val | tile187_jtag_ucb_val | tile203_jtag_ucb_val | tile219_jtag_ucb_val | tile235_jtag_ucb_val | tile251_jtag_ucb_val | tile12_jtag_ucb_val | tile28_jtag_ucb_val | tile44_jtag_ucb_val | tile60_jtag_ucb_val | tile76_jtag_ucb_val | tile92_jtag_ucb_val | tile108_jtag_ucb_val | tile124_jtag_ucb_val | tile140_jtag_ucb_val | tile156_jtag_ucb_val | tile172_jtag_ucb_val | tile188_jtag_ucb_val | tile204_jtag_ucb_val | tile220_jtag_ucb_val | tile236_jtag_ucb_val | tile252_jtag_ucb_val | tile13_jtag_ucb_val | tile29_jtag_ucb_val | tile45_jtag_ucb_val | tile61_jtag_ucb_val | tile77_jtag_ucb_val | tile93_jtag_ucb_val | tile109_jtag_ucb_val | tile125_jtag_ucb_val | tile141_jtag_ucb_val | tile157_jtag_ucb_val | tile173_jtag_ucb_val | tile189_jtag_ucb_val | tile205_jtag_ucb_val | tile221_jtag_ucb_val | tile237_jtag_ucb_val | tile253_jtag_ucb_val | tile14_jtag_ucb_val | tile30_jtag_ucb_val | tile46_jtag_ucb_val | tile62_jtag_ucb_val | tile78_jtag_ucb_val | tile94_jtag_ucb_val | tile110_jtag_ucb_val | tile126_jtag_ucb_val | tile142_jtag_ucb_val | tile158_jtag_ucb_val | tile174_jtag_ucb_val | tile190_jtag_ucb_val | tile206_jtag_ucb_val | tile222_jtag_ucb_val | tile238_jtag_ucb_val | tile254_jtag_ucb_val | tile15_jtag_ucb_val | tile31_jtag_ucb_val | tile47_jtag_ucb_val | tile63_jtag_ucb_val | tile79_jtag_ucb_val | tile95_jtag_ucb_val | tile111_jtag_ucb_val | tile127_jtag_ucb_val | tile143_jtag_ucb_val | tile159_jtag_ucb_val | tile175_jtag_ucb_val | tile191_jtag_ucb_val | tile207_jtag_ucb_val | tile223_jtag_ucb_val | tile239_jtag_ucb_val | tile255_jtag_ucb_val;
assign tiles_jtag_ucb_data = tile0_jtag_ucb_data | tile16_jtag_ucb_data | tile32_jtag_ucb_data | tile48_jtag_ucb_data | tile64_jtag_ucb_data | tile80_jtag_ucb_data | tile96_jtag_ucb_data | tile112_jtag_ucb_data | tile128_jtag_ucb_data | tile144_jtag_ucb_data | tile160_jtag_ucb_data | tile176_jtag_ucb_data | tile192_jtag_ucb_data | tile208_jtag_ucb_data | tile224_jtag_ucb_data | tile240_jtag_ucb_data | tile1_jtag_ucb_data | tile17_jtag_ucb_data | tile33_jtag_ucb_data | tile49_jtag_ucb_data | tile65_jtag_ucb_data | tile81_jtag_ucb_data | tile97_jtag_ucb_data | tile113_jtag_ucb_data | tile129_jtag_ucb_data | tile145_jtag_ucb_data | tile161_jtag_ucb_data | tile177_jtag_ucb_data | tile193_jtag_ucb_data | tile209_jtag_ucb_data | tile225_jtag_ucb_data | tile241_jtag_ucb_data | tile2_jtag_ucb_data | tile18_jtag_ucb_data | tile34_jtag_ucb_data | tile50_jtag_ucb_data | tile66_jtag_ucb_data | tile82_jtag_ucb_data | tile98_jtag_ucb_data | tile114_jtag_ucb_data | tile130_jtag_ucb_data | tile146_jtag_ucb_data | tile162_jtag_ucb_data | tile178_jtag_ucb_data | tile194_jtag_ucb_data | tile210_jtag_ucb_data | tile226_jtag_ucb_data | tile242_jtag_ucb_data | tile3_jtag_ucb_data | tile19_jtag_ucb_data | tile35_jtag_ucb_data | tile51_jtag_ucb_data | tile67_jtag_ucb_data | tile83_jtag_ucb_data | tile99_jtag_ucb_data | tile115_jtag_ucb_data | tile131_jtag_ucb_data | tile147_jtag_ucb_data | tile163_jtag_ucb_data | tile179_jtag_ucb_data | tile195_jtag_ucb_data | tile211_jtag_ucb_data | tile227_jtag_ucb_data | tile243_jtag_ucb_data | tile4_jtag_ucb_data | tile20_jtag_ucb_data | tile36_jtag_ucb_data | tile52_jtag_ucb_data | tile68_jtag_ucb_data | tile84_jtag_ucb_data | tile100_jtag_ucb_data | tile116_jtag_ucb_data | tile132_jtag_ucb_data | tile148_jtag_ucb_data | tile164_jtag_ucb_data | tile180_jtag_ucb_data | tile196_jtag_ucb_data | tile212_jtag_ucb_data | tile228_jtag_ucb_data | tile244_jtag_ucb_data | tile5_jtag_ucb_data | tile21_jtag_ucb_data | tile37_jtag_ucb_data | tile53_jtag_ucb_data | tile69_jtag_ucb_data | tile85_jtag_ucb_data | tile101_jtag_ucb_data | tile117_jtag_ucb_data | tile133_jtag_ucb_data | tile149_jtag_ucb_data | tile165_jtag_ucb_data | tile181_jtag_ucb_data | tile197_jtag_ucb_data | tile213_jtag_ucb_data | tile229_jtag_ucb_data | tile245_jtag_ucb_data | tile6_jtag_ucb_data | tile22_jtag_ucb_data | tile38_jtag_ucb_data | tile54_jtag_ucb_data | tile70_jtag_ucb_data | tile86_jtag_ucb_data | tile102_jtag_ucb_data | tile118_jtag_ucb_data | tile134_jtag_ucb_data | tile150_jtag_ucb_data | tile166_jtag_ucb_data | tile182_jtag_ucb_data | tile198_jtag_ucb_data | tile214_jtag_ucb_data | tile230_jtag_ucb_data | tile246_jtag_ucb_data | tile7_jtag_ucb_data | tile23_jtag_ucb_data | tile39_jtag_ucb_data | tile55_jtag_ucb_data | tile71_jtag_ucb_data | tile87_jtag_ucb_data | tile103_jtag_ucb_data | tile119_jtag_ucb_data | tile135_jtag_ucb_data | tile151_jtag_ucb_data | tile167_jtag_ucb_data | tile183_jtag_ucb_data | tile199_jtag_ucb_data | tile215_jtag_ucb_data | tile231_jtag_ucb_data | tile247_jtag_ucb_data | tile8_jtag_ucb_data | tile24_jtag_ucb_data | tile40_jtag_ucb_data | tile56_jtag_ucb_data | tile72_jtag_ucb_data | tile88_jtag_ucb_data | tile104_jtag_ucb_data | tile120_jtag_ucb_data | tile136_jtag_ucb_data | tile152_jtag_ucb_data | tile168_jtag_ucb_data | tile184_jtag_ucb_data | tile200_jtag_ucb_data | tile216_jtag_ucb_data | tile232_jtag_ucb_data | tile248_jtag_ucb_data | tile9_jtag_ucb_data | tile25_jtag_ucb_data | tile41_jtag_ucb_data | tile57_jtag_ucb_data | tile73_jtag_ucb_data | tile89_jtag_ucb_data | tile105_jtag_ucb_data | tile121_jtag_ucb_data | tile137_jtag_ucb_data | tile153_jtag_ucb_data | tile169_jtag_ucb_data | tile185_jtag_ucb_data | tile201_jtag_ucb_data | tile217_jtag_ucb_data | tile233_jtag_ucb_data | tile249_jtag_ucb_data | tile10_jtag_ucb_data | tile26_jtag_ucb_data | tile42_jtag_ucb_data | tile58_jtag_ucb_data | tile74_jtag_ucb_data | tile90_jtag_ucb_data | tile106_jtag_ucb_data | tile122_jtag_ucb_data | tile138_jtag_ucb_data | tile154_jtag_ucb_data | tile170_jtag_ucb_data | tile186_jtag_ucb_data | tile202_jtag_ucb_data | tile218_jtag_ucb_data | tile234_jtag_ucb_data | tile250_jtag_ucb_data | tile11_jtag_ucb_data | tile27_jtag_ucb_data | tile43_jtag_ucb_data | tile59_jtag_ucb_data | tile75_jtag_ucb_data | tile91_jtag_ucb_data | tile107_jtag_ucb_data | tile123_jtag_ucb_data | tile139_jtag_ucb_data | tile155_jtag_ucb_data | tile171_jtag_ucb_data | tile187_jtag_ucb_data | tile203_jtag_ucb_data | tile219_jtag_ucb_data | tile235_jtag_ucb_data | tile251_jtag_ucb_data | tile12_jtag_ucb_data | tile28_jtag_ucb_data | tile44_jtag_ucb_data | tile60_jtag_ucb_data | tile76_jtag_ucb_data | tile92_jtag_ucb_data | tile108_jtag_ucb_data | tile124_jtag_ucb_data | tile140_jtag_ucb_data | tile156_jtag_ucb_data | tile172_jtag_ucb_data | tile188_jtag_ucb_data | tile204_jtag_ucb_data | tile220_jtag_ucb_data | tile236_jtag_ucb_data | tile252_jtag_ucb_data | tile13_jtag_ucb_data | tile29_jtag_ucb_data | tile45_jtag_ucb_data | tile61_jtag_ucb_data | tile77_jtag_ucb_data | tile93_jtag_ucb_data | tile109_jtag_ucb_data | tile125_jtag_ucb_data | tile141_jtag_ucb_data | tile157_jtag_ucb_data | tile173_jtag_ucb_data | tile189_jtag_ucb_data | tile205_jtag_ucb_data | tile221_jtag_ucb_data | tile237_jtag_ucb_data | tile253_jtag_ucb_data | tile14_jtag_ucb_data | tile30_jtag_ucb_data | tile46_jtag_ucb_data | tile62_jtag_ucb_data | tile78_jtag_ucb_data | tile94_jtag_ucb_data | tile110_jtag_ucb_data | tile126_jtag_ucb_data | tile142_jtag_ucb_data | tile158_jtag_ucb_data | tile174_jtag_ucb_data | tile190_jtag_ucb_data | tile206_jtag_ucb_data | tile222_jtag_ucb_data | tile238_jtag_ucb_data | tile254_jtag_ucb_data | tile15_jtag_ucb_data | tile31_jtag_ucb_data | tile47_jtag_ucb_data | tile63_jtag_ucb_data | tile79_jtag_ucb_data | tile95_jtag_ucb_data | tile111_jtag_ucb_data | tile127_jtag_ucb_data | tile143_jtag_ucb_data | tile159_jtag_ucb_data | tile175_jtag_ucb_data | tile191_jtag_ucb_data | tile207_jtag_ucb_data | tile223_jtag_ucb_data | tile239_jtag_ucb_data | tile255_jtag_ucb_data;


   /////////////////////////
   // Sub-module Instances
   /////////////////////////

   // Need to generate clocks from MMCM for standalone chip FPGA synthesis
`ifdef PITON_FPGA_CLKS_GEN
   // Generate core_ref_clk
   clk_mmcm_chip clk_mmcm (
      .clk_in1_p(clk_osc_p),
      .clk_in1_n(clk_osc_n),

      .reset(1'b0),
      .locked(mmcm_locked),

      .core_ref_clk(core_ref_clk)
   );
`endif // endif PITON_FPGA_CLKS_GEN

`ifndef PITON_NO_CHIP_BRIDGE
`ifdef PITON_CHIP_FPGA
   // Generate io_clk from input
   IBUFGDS #(.DIFF_TERM("TRUE")) intf_chip_clk_ibufgds(
      .I(intf_chip_clk_p),
      .IB(intf_chip_clk_n),
      .O(io_clk)
   );
   // Output io_clk to intf
   OBUFDS chip_intf_clk_obufds(
      .I(io_clk),
      .O(chip_intf_clk_p),
      .OB(chip_intf_clk_n)
   );

   // Differential to single ended conversion for interface
   OBUFDS chip_intf_data_obufds[31:0] (
      .I(chip_intf_data),
      .O(chip_intf_data_p),
      .OB(chip_intf_data_n)
   );
   OBUFDS chip_intf_channel_obufds[1:0] (
      .I(chip_intf_channel),
      .O(chip_intf_channel_p),
      .OB(chip_intf_channel_n)
   );
   IBUFDS  #(.DIFF_TERM("TRUE")) chip_intf_credit_back_ibufds[2:0] (
      .I(chip_intf_credit_back_p),
      .IB(chip_intf_credit_back_n),
      .O(chip_intf_credit_back)
   );
   IBUFDS #(.DIFF_TERM("TRUE")) intf_chip_data_ibufds[31:0] (
      .I(intf_chip_data_p),
      .IB(intf_chip_data_n),
      .O(intf_chip_data)
   );
   IBUFDS #(.DIFF_TERM("TRUE")) intf_chip_channel_ibufds[1:0] (
      .I(intf_chip_channel_p),
      .IB(intf_chip_channel_n),
      .O(intf_chip_channel)
   );
   OBUFDS intf_chip_credit_back_obufds[2:0] (
      .I(intf_chip_credit_back),
      .O(intf_chip_credit_back_p),
      .OB(intf_chip_credit_back_n)
   );
`endif // endif PITON_CHIP_FPGA
`endif // endif PITON_NO_CHIP_BRIDGE

   // Off-Chip Interface Block

   OCI oci_inst (
   // Outside
   .slew                (slew),
   .impsel1                (impsel1),
   .impsel2                (impsel2),
   .core_ref_clk           (core_ref_clk),
   .io_clk                 (io_clk),
`ifndef PITON_CHIP_FPGA
   .rst_n                  (rst_n),
`else // ifndef PITON_CHIP_FPGA
   .rst_n                       (rst_n & (~chipset_prsnt_n)),
`endif
   .pll_rst_n              (pll_rst_n),
   .pll_rangea             (pll_rangea),
   .clk_mux_sel               (clk_mux_sel),
   .clk_en                 (clk_en),
   .pll_bypass             (pll_bypass),
   .async_mux              (async_mux),
   .oram_on                (oram_on),
   .oram_traffic_gen       (oram_traffic_gen),
   .oram_dummy_gen            (oram_dummy_gen),
   .pll_lock               (pll_lock),
   .jtag_clk               (jtag_clk),
   .jtag_rst_l             (jtag_rst_l),
   .jtag_modesel           (jtag_modesel),
   .jtag_datain               (jtag_datain),
   .jtag_dataout           (jtag_dataout),
`ifndef PITON_NO_CHIP_BRIDGE
   .intf_chip_data            (intf_chip_data),
   .intf_chip_channel         (intf_chip_channel),
   .intf_chip_credit_back     (intf_chip_credit_back),
   .chip_intf_data            (chip_intf_data),
   .chip_intf_channel         (chip_intf_channel),
   .chip_intf_credit_back     (chip_intf_credit_back),
`else // ifdef PITON_NO_CHIP_BRIDGE
   .intf_chip_data              (),
   .intf_chip_channel           (),
   .intf_chip_credit_back       (),
   .chip_intf_data              (),
   .chip_intf_channel           (),
   .chip_intf_credit_back       (),
`endif // endif PITON_NO_CHIP_BRIDGE
   // Inside
   .core_ref_clk_inter        (core_ref_clk_inter),
   .io_clk_inter           (io_clk_inter),
   .rst_n_inter               (rst_n_inter),
   .pll_rst_n_inter           (pll_rst_n_inter),
   .pll_rangea_inter       (pll_rangea_inter),
   .clk_mux_sel_inter         (clk_mux_sel_inter),
   .clk_en_inter           (clk_en_inter),
   .pll_bypass_inter       (pll_bypass_inter),
   .async_mux_inter           (async_mux_inter),
   .oram_on_inter          (oram_on_inter),
   .oram_traffic_gen_inter    (oram_traffic_gen_inter),
   .oram_dummy_gen_inter      (oram_dummy_gen_inter),
   .pll_lock_inter            (pll_lock_inter),
   .jtag_clk_inter            (jtag_clk_inter),
   .jtag_rst_l_inter       (jtag_rst_l_inter),
   .jtag_modesel_inter        (jtag_modesel_inter),
   .jtag_datain_inter         (jtag_datain_inter),
   .jtag_dataout_inter        (jtag_dataout_inter),
   .intf_chip_data_inter      (intf_chip_data_inter),
   .intf_chip_channel_inter      (intf_chip_channel_inter),
   .intf_chip_credit_back_inter  (intf_chip_credit_back_inter),
   .chip_intf_data_inter      (chip_intf_data_inter),
   .chip_intf_channel_inter      (chip_intf_channel_inter),
   .chip_intf_credit_back_inter  (chip_intf_credit_back_inter) );

   // PLL and clock mux.  See above for alternatives
   clk_se_to_diff ref_clk_converter (
       .clk_se  (core_ref_clk_inter),
       .clk_p   (core_ref_clk_inter_t),
       .clk_n   (core_ref_clk_inter_c)
   );
   clk_mux clock_mux (
       .clk0_p(core_ref_clk_inter_t),
       .clk0_n(core_ref_clk_inter_c),
       .clk1_p(1'b1),
       .clk1_n(1'b0),
       .clk2(pll_clk),

       .sel(clk_mux_sel_inter),

       .clk_muxed(clk_muxed)
   );
   pll_top pll_top (
      .clk_locked(pll_lock_inter),
      .clk_out(pll_clk),

      .rangeA(pll_rangea_inter),
      .bypass_en(pll_bypass_inter),
      .ref_clk(core_ref_clk_inter),
      .rst(~pll_rst_n_inter)
   );

   // reset synchronizer, might need to be placed near the
   //   pll or clock source so that reset signal has the same propagation
   //   as clock for better timing
   // materials on reset tree and placement
   // http://www.sunburst-design.com/papers/CummingsSNUG2002SJ_Resets.pdf
   synchronizer rst_sync (
      .clk(clk_muxed),
      .presyncdata(rst_n_inter),
      .syncdata(rst_n_inter_sync)
   );
   synchronizer io_clk_rst_sync (
      .clk(io_clk_inter),
      .presyncdata(rst_n_inter),
      .syncdata(io_clk_rst_n_inter_sync)
   );
   synchronizer jtag_rst_sync (
      .clk(clk_muxed),
      .presyncdata(jtag_rst_l_inter),
      .syncdata(jtag_rst_l_inter_sync)
   );

`ifndef PITON_NO_CHIP_BRIDGE
   // Chip to FPGA bridge
   chip_bridge chip_intf(
       // Xilinx afifos want asynchronous reset, so need to passs that in
       // and do internal synchronizeation
`ifdef PITON_PROTO
       .rst_n                  (rst_n_inter),
`else // ifndef PITON_FPGA_SYNTH
       .rst_n                  (rst_n_inter_sync_f),
`endif
       .chip_clk               (clk_muxed),
       .intcnct_clk            (io_clk_inter),
       .async_mux              (async_mux_inter),
       .network_out_1          (chip_intf_noc1_data),
       .network_out_2          (chip_intf_noc2_data),
       .network_out_3          (chip_intf_noc3_data),
       .data_out_val_1         (chip_intf_noc1_valid),
       .data_out_val_2         (chip_intf_noc2_valid),
       .data_out_val_3         (chip_intf_noc3_valid),
       .data_out_rdy_1         (chip_intf_noc1_rdy),
       .data_out_rdy_2         (chip_intf_noc2_rdy),
       .data_out_rdy_3         (chip_intf_noc3_rdy),
       .intcnct_data_in        (intf_chip_data_inter_buf_f),
       .intcnct_channel_in     (intf_chip_channel_inter_buf_f),
       .intcnct_credit_back_in (intf_chip_credit_back_inter),
       .network_in_1           (intf_chip_noc1_data),
       .network_in_2           (intf_chip_noc2_data),
       .network_in_3           (intf_chip_noc3_data),
       .data_in_val_1          (intf_chip_noc1_valid),
       .data_in_val_2          (intf_chip_noc2_valid),
       .data_in_val_3          (intf_chip_noc3_valid),
       .data_in_rdy_1          (intf_chip_noc1_rdy),
       .data_in_rdy_2          (intf_chip_noc2_rdy),
       .data_in_rdy_3          (intf_chip_noc3_rdy),
       .intcnct_data_out       (chip_intf_data_inter),
       .intcnct_channel_out    (chip_intf_channel_inter),
       .intcnct_credit_back_out(chip_intf_credit_back_inter_buf_f)
   );

   // Chip Bridge val/rdy to credit

   valrdy_to_credit #(4, 3) chip_from_intf_noc1_v2c(
      .clk(clk_muxed),
      .reset(~rst_n_inter_sync_f),
      .data_in(intf_chip_noc1_data),
      .valid_in(intf_chip_noc1_valid),
      .ready_in(intf_chip_noc1_rdy),

      .data_out(offchip_processor_noc1_data),           // Data
      .valid_out(offchip_processor_noc1_valid),       // Val signal
      .yummy_out(offchip_processor_noc1_yummy)    // Yummy signal
   );

   credit_to_valrdy chip_to_intf_noc1_c2v(
      .clk(clk_muxed),
      .reset(~rst_n_inter_sync_f),
      .data_in(processor_offchip_noc1_data),
      .valid_in(processor_offchip_noc1_valid),
      .yummy_in(processor_offchip_noc1_yummy),

      .data_out(chip_intf_noc1_data),           // Data
      .valid_out(chip_intf_noc1_valid),       // Val signal from dynamic network to processor
      .ready_out(chip_intf_noc1_rdy)    // Rdy signal from processor to dynamic network
   );

   valrdy_to_credit #(4, 3) chip_from_intf_noc2_v2c(
      .clk(clk_muxed),
      .reset(~rst_n_inter_sync_f),
      .data_in(intf_chip_noc2_data),
      .valid_in(intf_chip_noc2_valid),
      .ready_in(intf_chip_noc2_rdy),

      .data_out(offchip_processor_noc2_data),           // Data
      .valid_out(offchip_processor_noc2_valid),       // Val signal
      .yummy_out(offchip_processor_noc2_yummy)    // Yummy signal
   );

   credit_to_valrdy chip_to_intf_noc2_c2v(
      .clk(clk_muxed),
      .reset(~rst_n_inter_sync_f),
      .data_in(processor_offchip_noc2_data),
      .valid_in(processor_offchip_noc2_valid),
      .yummy_in(processor_offchip_noc2_yummy),

      .data_out(chip_intf_noc2_data),           // Data
      .valid_out(chip_intf_noc2_valid),       // Val signal from dynamic network to processor
      .ready_out(chip_intf_noc2_rdy)    // Rdy signal from processor to dynamic network
   );

   valrdy_to_credit #(4, 3) chip_from_intf_noc3_v2c(
      .clk(clk_muxed),
      .reset(~rst_n_inter_sync_f),
      .data_in(intf_chip_noc3_data),
      .valid_in(intf_chip_noc3_valid),
      .ready_in(intf_chip_noc3_rdy),

      .data_out(offchip_processor_noc3_data),           // Data
      .valid_out(offchip_processor_noc3_valid),       // Val signal
      .yummy_out(offchip_processor_noc3_yummy)    // Yummy signal
   );

   credit_to_valrdy chip_to_intf_noc3_c2v(
      .clk(clk_muxed),
      .reset(~rst_n_inter_sync_f),
      .data_in(processor_offchip_noc3_data),
      .valid_in(processor_offchip_noc3_valid),
      .yummy_in(processor_offchip_noc3_yummy),

      .data_out(chip_intf_noc3_data),           // Data
      .valid_out(chip_intf_noc3_valid),       // Val signal from dynamic network to processor
      .ready_out(chip_intf_noc3_rdy)    // Rdy signal from processor to dynamic network
   );
`endif // endif PITON_NO_CHIP_BRIDGE

`ifdef ORAM_ON
   oram_top oram_top(
      .clk(clk_muxed),
      .rst_n(rst_n_inter_sync),
      .clk_en(ctap_oram_clk_en && clk_en_inter),
      .oram_on(oram_on_inter),
      .oram_traffic_gen(oram_traffic_gen_inter),
      .oram_dummy_gen(oram_dummy_gen_inter),

      //from noc2
      .proc_oram_valid(proc_oram_valid),
      .proc_oram_data(proc_oram_data),
      .proc_oram_yummy(proc_oram_yummy_oram),

      //to noc3
      .oram_proc_valid(oram_proc_valid_oram),
      .oram_proc_data(oram_proc_data_oram),
      .oram_proc_yummy(oram_proc_yummy),

      //from noc3
      .offchip_oram_valid(offchip_oram_valid),
      .offchip_oram_data(offchip_oram_data),
      .offchip_oram_yummy(offchip_oram_yummy_oram),

      //to noc2
      .oram_offchip_valid(oram_offchip_valid_oram),
      .oram_offchip_data(oram_offchip_data_oram),
      .oram_offchip_yummy(oram_offchip_yummy),

      // oram-jtag
      .ctap_oram_req_val(ctap_oram_req_val),
      // .ctap_oram_req_misc(ctap_oram_req_misc),
      .oram_ctap_res_data(oram_ctap_res_data)
      // .ctap_oram_bist_command(ctap_oram_bist_command),
      // .ctap_oram_bist_data(ctap_oram_bist_data),
      // .oram_ctap_sram_data(oram_ctap_sram_data)
   );
`endif // endif ORAM_ON

   // on-chip jtag interface & test access port
   jtag jtag_port(
      .clk(clk_muxed),
      .rst_n(rst_n_inter_sync_f),
      .jtag_clk(jtag_clk_inter),
      .jtag_rst_l(jtag_rst_l_inter_sync),
      .jtag_modesel(jtag_modesel_inter),
      .jtag_datain(jtag_datain_inter),
      .jtag_dataout(jtag_dataout_inter),
      .jtag_dataout_en(),
      .jtag_tiles_ucb_val(jtag_tiles_ucb_val),
      .jtag_tiles_ucb_data(jtag_tiles_ucb_data),
      .tiles_jtag_ucb_val(tiles_jtag_ucb_val),
      .tiles_jtag_ucb_data(tiles_jtag_ucb_data),

      .ctap_oram_req_val(ctap_oram_req_val),
      .ctap_oram_req_misc(ctap_oram_req_misc),
      .oram_ctap_res_data(oram_ctap_res_data),
      // .ctap_oram_bist_command(ctap_oram_bist_command),
      // .ctap_oram_bist_data(ctap_oram_bist_data),
      // .oram_ctap_sram_data(oram_ctap_sram_data),

      .ctap_clk_en(ctap_clk_en_inter),
      .ctap_oram_clk_en(ctap_oram_clk_en)
   );

   // generate the cross bars


    wire [31:0] default_total_num_tiles;
    assign default_total_num_tiles = `PITON_NUM_TILES;
    // Generate tile instances

tile
tile0 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[0] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd0),
    .default_coreid_y           (8'd0),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd0)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[0]   )
    ,.unavailable_o       ( unavailable_o[0] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[0]   )
    ,.ipi_i               ( ipi_i[0]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[0*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile0_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile0_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( dummy_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_0_1_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( offchip_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_1_0_out_N_noc1_data   ),
    .dyn0_validIn_N      ( dummy_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_0_1_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( offchip_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_1_0_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( dummy_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_0_1_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( offchip_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_1_0_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_0_0_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_0_0_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_0_0_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_0_0_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_0_0_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_0_0_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_0_0_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_0_0_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_0_0_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_0_0_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_0_0_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_0_0_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( dummy_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_0_1_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( offchip_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_1_0_out_N_noc2_data   ),
    .dyn1_validIn_N      ( dummy_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_0_1_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( offchip_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_1_0_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( dummy_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_0_1_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( offchip_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_1_0_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_0_0_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_0_0_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_0_0_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_0_0_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_0_0_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_0_0_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_0_0_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_0_0_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_0_0_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_0_0_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_0_0_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_0_0_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( dummy_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_0_1_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( offchip_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_1_0_out_N_noc3_data   ),
    .dyn2_validIn_N      ( dummy_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_0_1_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( offchip_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_1_0_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( dummy_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_0_1_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( offchip_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_1_0_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_0_0_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_0_0_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_0_0_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_0_0_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_0_0_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_0_0_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_0_0_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_0_0_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_0_0_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_0_0_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_0_0_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_0_0_out_S_noc3_yummy )
);


tile
tile16 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[16] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd0),
    .default_coreid_y           (8'd1),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd16)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[16]   )
    ,.unavailable_o       ( unavailable_o[16] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[16]   )
    ,.ipi_i               ( ipi_i[16]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[16*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile16_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile16_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_0_0_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_1_1_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( dummy_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_2_0_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_0_0_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_1_1_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( dummy_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_2_0_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_0_0_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_1_1_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( dummy_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_2_0_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_1_0_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_1_0_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_1_0_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_1_0_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_1_0_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_1_0_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_1_0_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_1_0_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_1_0_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_1_0_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_1_0_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_1_0_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_0_0_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_1_1_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( dummy_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_2_0_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_0_0_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_1_1_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( dummy_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_2_0_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_0_0_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_1_1_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( dummy_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_2_0_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_1_0_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_1_0_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_1_0_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_1_0_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_1_0_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_1_0_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_1_0_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_1_0_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_1_0_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_1_0_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_1_0_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_1_0_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_0_0_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_1_1_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( dummy_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_2_0_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_0_0_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_1_1_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( dummy_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_2_0_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_0_0_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_1_1_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( dummy_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_2_0_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_1_0_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_1_0_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_1_0_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_1_0_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_1_0_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_1_0_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_1_0_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_1_0_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_1_0_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_1_0_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_1_0_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_1_0_out_S_noc3_yummy )
);


tile
tile32 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[32] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd0),
    .default_coreid_y           (8'd2),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd32)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[32]   )
    ,.unavailable_o       ( unavailable_o[32] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[32]   )
    ,.ipi_i               ( ipi_i[32]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[32*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile32_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile32_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_1_0_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_2_1_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( dummy_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_3_0_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_1_0_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_2_1_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( dummy_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_3_0_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_1_0_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_2_1_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( dummy_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_3_0_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_2_0_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_2_0_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_2_0_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_2_0_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_2_0_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_2_0_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_2_0_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_2_0_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_2_0_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_2_0_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_2_0_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_2_0_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_1_0_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_2_1_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( dummy_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_3_0_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_1_0_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_2_1_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( dummy_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_3_0_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_1_0_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_2_1_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( dummy_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_3_0_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_2_0_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_2_0_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_2_0_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_2_0_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_2_0_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_2_0_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_2_0_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_2_0_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_2_0_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_2_0_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_2_0_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_2_0_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_1_0_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_2_1_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( dummy_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_3_0_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_1_0_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_2_1_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( dummy_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_3_0_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_1_0_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_2_1_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( dummy_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_3_0_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_2_0_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_2_0_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_2_0_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_2_0_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_2_0_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_2_0_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_2_0_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_2_0_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_2_0_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_2_0_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_2_0_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_2_0_out_S_noc3_yummy )
);


tile
tile48 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[48] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd0),
    .default_coreid_y           (8'd3),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd48)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[48]   )
    ,.unavailable_o       ( unavailable_o[48] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[48]   )
    ,.ipi_i               ( ipi_i[48]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[48*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile48_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile48_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_2_0_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_3_1_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( dummy_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_4_0_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_2_0_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_3_1_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( dummy_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_4_0_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_2_0_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_3_1_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( dummy_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_4_0_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_3_0_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_3_0_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_3_0_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_3_0_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_3_0_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_3_0_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_3_0_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_3_0_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_3_0_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_3_0_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_3_0_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_3_0_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_2_0_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_3_1_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( dummy_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_4_0_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_2_0_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_3_1_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( dummy_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_4_0_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_2_0_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_3_1_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( dummy_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_4_0_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_3_0_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_3_0_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_3_0_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_3_0_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_3_0_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_3_0_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_3_0_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_3_0_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_3_0_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_3_0_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_3_0_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_3_0_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_2_0_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_3_1_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( dummy_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_4_0_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_2_0_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_3_1_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( dummy_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_4_0_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_2_0_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_3_1_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( dummy_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_4_0_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_3_0_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_3_0_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_3_0_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_3_0_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_3_0_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_3_0_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_3_0_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_3_0_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_3_0_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_3_0_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_3_0_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_3_0_out_S_noc3_yummy )
);


tile
tile64 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[64] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd0),
    .default_coreid_y           (8'd4),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd64)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[64]   )
    ,.unavailable_o       ( unavailable_o[64] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[64]   )
    ,.ipi_i               ( ipi_i[64]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[64*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile64_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile64_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_3_0_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_4_1_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( dummy_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_5_0_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_3_0_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_4_1_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( dummy_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_5_0_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_3_0_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_4_1_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( dummy_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_5_0_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_4_0_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_4_0_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_4_0_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_4_0_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_4_0_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_4_0_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_4_0_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_4_0_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_4_0_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_4_0_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_4_0_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_4_0_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_3_0_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_4_1_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( dummy_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_5_0_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_3_0_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_4_1_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( dummy_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_5_0_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_3_0_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_4_1_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( dummy_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_5_0_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_4_0_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_4_0_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_4_0_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_4_0_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_4_0_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_4_0_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_4_0_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_4_0_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_4_0_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_4_0_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_4_0_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_4_0_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_3_0_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_4_1_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( dummy_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_5_0_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_3_0_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_4_1_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( dummy_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_5_0_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_3_0_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_4_1_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( dummy_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_5_0_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_4_0_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_4_0_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_4_0_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_4_0_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_4_0_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_4_0_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_4_0_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_4_0_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_4_0_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_4_0_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_4_0_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_4_0_out_S_noc3_yummy )
);


tile
tile80 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[80] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd0),
    .default_coreid_y           (8'd5),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd80)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[80]   )
    ,.unavailable_o       ( unavailable_o[80] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[80]   )
    ,.ipi_i               ( ipi_i[80]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[80*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile80_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile80_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_4_0_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_5_1_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( dummy_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_6_0_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_4_0_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_5_1_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( dummy_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_6_0_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_4_0_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_5_1_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( dummy_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_6_0_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_5_0_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_5_0_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_5_0_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_5_0_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_5_0_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_5_0_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_5_0_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_5_0_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_5_0_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_5_0_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_5_0_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_5_0_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_4_0_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_5_1_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( dummy_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_6_0_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_4_0_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_5_1_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( dummy_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_6_0_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_4_0_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_5_1_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( dummy_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_6_0_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_5_0_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_5_0_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_5_0_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_5_0_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_5_0_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_5_0_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_5_0_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_5_0_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_5_0_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_5_0_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_5_0_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_5_0_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_4_0_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_5_1_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( dummy_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_6_0_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_4_0_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_5_1_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( dummy_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_6_0_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_4_0_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_5_1_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( dummy_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_6_0_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_5_0_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_5_0_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_5_0_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_5_0_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_5_0_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_5_0_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_5_0_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_5_0_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_5_0_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_5_0_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_5_0_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_5_0_out_S_noc3_yummy )
);


tile
tile96 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[96] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd0),
    .default_coreid_y           (8'd6),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd96)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[96]   )
    ,.unavailable_o       ( unavailable_o[96] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[96]   )
    ,.ipi_i               ( ipi_i[96]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[96*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile96_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile96_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_5_0_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_6_1_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( dummy_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_7_0_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_5_0_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_6_1_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( dummy_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_7_0_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_5_0_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_6_1_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( dummy_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_7_0_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_6_0_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_6_0_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_6_0_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_6_0_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_6_0_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_6_0_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_6_0_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_6_0_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_6_0_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_6_0_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_6_0_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_6_0_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_5_0_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_6_1_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( dummy_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_7_0_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_5_0_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_6_1_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( dummy_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_7_0_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_5_0_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_6_1_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( dummy_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_7_0_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_6_0_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_6_0_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_6_0_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_6_0_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_6_0_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_6_0_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_6_0_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_6_0_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_6_0_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_6_0_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_6_0_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_6_0_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_5_0_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_6_1_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( dummy_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_7_0_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_5_0_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_6_1_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( dummy_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_7_0_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_5_0_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_6_1_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( dummy_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_7_0_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_6_0_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_6_0_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_6_0_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_6_0_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_6_0_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_6_0_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_6_0_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_6_0_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_6_0_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_6_0_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_6_0_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_6_0_out_S_noc3_yummy )
);


tile
tile112 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[112] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd0),
    .default_coreid_y           (8'd7),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd112)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[112]   )
    ,.unavailable_o       ( unavailable_o[112] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[112]   )
    ,.ipi_i               ( ipi_i[112]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[112*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile112_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile112_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_6_0_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_7_1_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( dummy_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_8_0_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_6_0_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_7_1_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( dummy_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_8_0_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_6_0_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_7_1_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( dummy_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_8_0_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_7_0_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_7_0_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_7_0_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_7_0_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_7_0_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_7_0_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_7_0_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_7_0_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_7_0_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_7_0_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_7_0_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_7_0_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_6_0_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_7_1_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( dummy_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_8_0_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_6_0_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_7_1_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( dummy_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_8_0_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_6_0_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_7_1_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( dummy_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_8_0_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_7_0_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_7_0_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_7_0_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_7_0_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_7_0_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_7_0_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_7_0_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_7_0_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_7_0_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_7_0_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_7_0_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_7_0_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_6_0_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_7_1_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( dummy_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_8_0_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_6_0_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_7_1_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( dummy_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_8_0_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_6_0_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_7_1_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( dummy_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_8_0_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_7_0_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_7_0_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_7_0_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_7_0_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_7_0_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_7_0_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_7_0_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_7_0_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_7_0_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_7_0_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_7_0_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_7_0_out_S_noc3_yummy )
);


tile
tile128 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[128] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd0),
    .default_coreid_y           (8'd8),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd128)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[128]   )
    ,.unavailable_o       ( unavailable_o[128] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[128]   )
    ,.ipi_i               ( ipi_i[128]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[128*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile128_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile128_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_7_0_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_8_1_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( dummy_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_9_0_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_7_0_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_8_1_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( dummy_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_9_0_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_7_0_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_8_1_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( dummy_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_9_0_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_8_0_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_8_0_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_8_0_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_8_0_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_8_0_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_8_0_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_8_0_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_8_0_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_8_0_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_8_0_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_8_0_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_8_0_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_7_0_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_8_1_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( dummy_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_9_0_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_7_0_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_8_1_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( dummy_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_9_0_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_7_0_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_8_1_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( dummy_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_9_0_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_8_0_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_8_0_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_8_0_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_8_0_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_8_0_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_8_0_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_8_0_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_8_0_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_8_0_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_8_0_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_8_0_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_8_0_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_7_0_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_8_1_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( dummy_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_9_0_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_7_0_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_8_1_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( dummy_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_9_0_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_7_0_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_8_1_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( dummy_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_9_0_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_8_0_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_8_0_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_8_0_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_8_0_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_8_0_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_8_0_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_8_0_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_8_0_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_8_0_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_8_0_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_8_0_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_8_0_out_S_noc3_yummy )
);


tile
tile144 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[144] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd0),
    .default_coreid_y           (8'd9),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd144)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[144]   )
    ,.unavailable_o       ( unavailable_o[144] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[144]   )
    ,.ipi_i               ( ipi_i[144]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[144*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile144_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile144_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_8_0_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_9_1_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( dummy_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_10_0_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_8_0_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_9_1_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( dummy_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_10_0_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_8_0_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_9_1_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( dummy_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_10_0_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_9_0_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_9_0_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_9_0_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_9_0_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_9_0_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_9_0_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_9_0_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_9_0_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_9_0_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_9_0_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_9_0_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_9_0_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_8_0_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_9_1_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( dummy_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_10_0_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_8_0_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_9_1_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( dummy_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_10_0_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_8_0_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_9_1_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( dummy_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_10_0_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_9_0_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_9_0_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_9_0_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_9_0_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_9_0_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_9_0_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_9_0_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_9_0_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_9_0_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_9_0_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_9_0_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_9_0_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_8_0_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_9_1_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( dummy_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_10_0_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_8_0_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_9_1_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( dummy_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_10_0_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_8_0_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_9_1_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( dummy_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_10_0_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_9_0_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_9_0_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_9_0_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_9_0_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_9_0_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_9_0_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_9_0_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_9_0_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_9_0_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_9_0_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_9_0_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_9_0_out_S_noc3_yummy )
);


tile
tile160 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[160] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd0),
    .default_coreid_y           (8'd10),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd160)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[160]   )
    ,.unavailable_o       ( unavailable_o[160] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[160]   )
    ,.ipi_i               ( ipi_i[160]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[160*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile160_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile160_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_9_0_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_10_1_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( dummy_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_11_0_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_9_0_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_10_1_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( dummy_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_11_0_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_9_0_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_10_1_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( dummy_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_11_0_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_10_0_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_10_0_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_10_0_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_10_0_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_10_0_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_10_0_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_10_0_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_10_0_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_10_0_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_10_0_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_10_0_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_10_0_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_9_0_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_10_1_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( dummy_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_11_0_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_9_0_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_10_1_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( dummy_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_11_0_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_9_0_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_10_1_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( dummy_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_11_0_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_10_0_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_10_0_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_10_0_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_10_0_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_10_0_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_10_0_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_10_0_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_10_0_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_10_0_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_10_0_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_10_0_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_10_0_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_9_0_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_10_1_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( dummy_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_11_0_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_9_0_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_10_1_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( dummy_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_11_0_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_9_0_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_10_1_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( dummy_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_11_0_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_10_0_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_10_0_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_10_0_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_10_0_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_10_0_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_10_0_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_10_0_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_10_0_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_10_0_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_10_0_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_10_0_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_10_0_out_S_noc3_yummy )
);


tile
tile176 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[176] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd0),
    .default_coreid_y           (8'd11),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd176)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[176]   )
    ,.unavailable_o       ( unavailable_o[176] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[176]   )
    ,.ipi_i               ( ipi_i[176]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[176*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile176_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile176_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_10_0_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_11_1_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( dummy_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_12_0_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_10_0_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_11_1_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( dummy_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_12_0_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_10_0_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_11_1_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( dummy_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_12_0_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_11_0_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_11_0_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_11_0_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_11_0_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_11_0_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_11_0_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_11_0_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_11_0_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_11_0_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_11_0_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_11_0_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_11_0_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_10_0_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_11_1_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( dummy_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_12_0_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_10_0_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_11_1_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( dummy_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_12_0_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_10_0_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_11_1_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( dummy_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_12_0_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_11_0_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_11_0_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_11_0_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_11_0_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_11_0_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_11_0_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_11_0_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_11_0_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_11_0_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_11_0_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_11_0_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_11_0_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_10_0_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_11_1_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( dummy_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_12_0_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_10_0_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_11_1_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( dummy_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_12_0_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_10_0_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_11_1_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( dummy_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_12_0_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_11_0_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_11_0_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_11_0_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_11_0_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_11_0_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_11_0_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_11_0_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_11_0_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_11_0_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_11_0_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_11_0_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_11_0_out_S_noc3_yummy )
);


tile
tile192 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[192] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd0),
    .default_coreid_y           (8'd12),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd192)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[192]   )
    ,.unavailable_o       ( unavailable_o[192] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[192]   )
    ,.ipi_i               ( ipi_i[192]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[192*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile192_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile192_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_11_0_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_12_1_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( dummy_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_13_0_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_11_0_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_12_1_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( dummy_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_13_0_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_11_0_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_12_1_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( dummy_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_13_0_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_12_0_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_12_0_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_12_0_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_12_0_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_12_0_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_12_0_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_12_0_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_12_0_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_12_0_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_12_0_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_12_0_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_12_0_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_11_0_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_12_1_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( dummy_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_13_0_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_11_0_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_12_1_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( dummy_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_13_0_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_11_0_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_12_1_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( dummy_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_13_0_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_12_0_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_12_0_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_12_0_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_12_0_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_12_0_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_12_0_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_12_0_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_12_0_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_12_0_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_12_0_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_12_0_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_12_0_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_11_0_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_12_1_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( dummy_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_13_0_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_11_0_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_12_1_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( dummy_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_13_0_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_11_0_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_12_1_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( dummy_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_13_0_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_12_0_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_12_0_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_12_0_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_12_0_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_12_0_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_12_0_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_12_0_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_12_0_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_12_0_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_12_0_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_12_0_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_12_0_out_S_noc3_yummy )
);


tile
tile208 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[208] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd0),
    .default_coreid_y           (8'd13),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd208)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[208]   )
    ,.unavailable_o       ( unavailable_o[208] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[208]   )
    ,.ipi_i               ( ipi_i[208]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[208*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile208_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile208_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_12_0_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_13_1_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( dummy_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_14_0_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_12_0_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_13_1_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( dummy_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_14_0_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_12_0_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_13_1_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( dummy_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_14_0_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_13_0_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_13_0_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_13_0_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_13_0_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_13_0_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_13_0_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_13_0_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_13_0_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_13_0_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_13_0_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_13_0_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_13_0_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_12_0_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_13_1_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( dummy_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_14_0_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_12_0_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_13_1_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( dummy_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_14_0_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_12_0_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_13_1_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( dummy_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_14_0_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_13_0_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_13_0_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_13_0_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_13_0_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_13_0_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_13_0_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_13_0_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_13_0_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_13_0_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_13_0_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_13_0_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_13_0_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_12_0_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_13_1_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( dummy_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_14_0_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_12_0_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_13_1_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( dummy_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_14_0_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_12_0_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_13_1_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( dummy_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_14_0_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_13_0_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_13_0_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_13_0_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_13_0_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_13_0_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_13_0_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_13_0_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_13_0_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_13_0_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_13_0_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_13_0_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_13_0_out_S_noc3_yummy )
);


tile
tile224 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[224] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd0),
    .default_coreid_y           (8'd14),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd224)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[224]   )
    ,.unavailable_o       ( unavailable_o[224] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[224]   )
    ,.ipi_i               ( ipi_i[224]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[224*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile224_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile224_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_13_0_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_14_1_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( dummy_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_15_0_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_13_0_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_14_1_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( dummy_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_15_0_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_13_0_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_14_1_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( dummy_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_15_0_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_14_0_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_14_0_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_14_0_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_14_0_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_14_0_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_14_0_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_14_0_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_14_0_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_14_0_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_14_0_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_14_0_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_14_0_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_13_0_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_14_1_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( dummy_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_15_0_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_13_0_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_14_1_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( dummy_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_15_0_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_13_0_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_14_1_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( dummy_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_15_0_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_14_0_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_14_0_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_14_0_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_14_0_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_14_0_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_14_0_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_14_0_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_14_0_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_14_0_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_14_0_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_14_0_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_14_0_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_13_0_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_14_1_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( dummy_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_15_0_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_13_0_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_14_1_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( dummy_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_15_0_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_13_0_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_14_1_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( dummy_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_15_0_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_14_0_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_14_0_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_14_0_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_14_0_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_14_0_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_14_0_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_14_0_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_14_0_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_14_0_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_14_0_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_14_0_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_14_0_out_S_noc3_yummy )
);


tile
tile240 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[240] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd0),
    .default_coreid_y           (8'd15),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd240)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[240]   )
    ,.unavailable_o       ( unavailable_o[240] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[240]   )
    ,.ipi_i               ( ipi_i[240]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[240*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile240_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile240_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_14_0_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_15_1_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( dummy_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( dummy_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_14_0_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_15_1_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( dummy_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( dummy_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_14_0_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_15_1_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( dummy_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( dummy_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_15_0_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_15_0_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_15_0_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_15_0_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_15_0_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_15_0_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_15_0_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_15_0_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_15_0_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_15_0_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_15_0_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_15_0_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_14_0_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_15_1_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( dummy_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( dummy_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_14_0_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_15_1_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( dummy_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( dummy_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_14_0_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_15_1_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( dummy_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( dummy_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_15_0_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_15_0_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_15_0_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_15_0_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_15_0_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_15_0_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_15_0_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_15_0_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_15_0_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_15_0_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_15_0_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_15_0_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_14_0_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_15_1_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( dummy_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( dummy_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_14_0_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_15_1_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( dummy_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( dummy_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_14_0_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_15_1_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( dummy_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( dummy_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_15_0_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_15_0_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_15_0_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_15_0_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_15_0_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_15_0_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_15_0_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_15_0_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_15_0_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_15_0_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_15_0_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_15_0_out_S_noc3_yummy )
);


tile
tile1 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[1] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd1),
    .default_coreid_y           (8'd0),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd1)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[1]   )
    ,.unavailable_o       ( unavailable_o[1] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[1]   )
    ,.ipi_i               ( ipi_i[1]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[1*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile1_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile1_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( dummy_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_0_2_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_0_0_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_1_1_out_N_noc1_data   ),
    .dyn0_validIn_N      ( dummy_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_0_2_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_0_0_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_1_1_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( dummy_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_0_2_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_0_0_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_1_1_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_0_1_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_0_1_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_0_1_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_0_1_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_0_1_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_0_1_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_0_1_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_0_1_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_0_1_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_0_1_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_0_1_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_0_1_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( dummy_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_0_2_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_0_0_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_1_1_out_N_noc2_data   ),
    .dyn1_validIn_N      ( dummy_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_0_2_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_0_0_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_1_1_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( dummy_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_0_2_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_0_0_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_1_1_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_0_1_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_0_1_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_0_1_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_0_1_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_0_1_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_0_1_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_0_1_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_0_1_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_0_1_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_0_1_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_0_1_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_0_1_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( dummy_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_0_2_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_0_0_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_1_1_out_N_noc3_data   ),
    .dyn2_validIn_N      ( dummy_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_0_2_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_0_0_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_1_1_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( dummy_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_0_2_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_0_0_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_1_1_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_0_1_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_0_1_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_0_1_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_0_1_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_0_1_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_0_1_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_0_1_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_0_1_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_0_1_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_0_1_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_0_1_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_0_1_out_S_noc3_yummy )
);


tile
tile17 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[17] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd1),
    .default_coreid_y           (8'd1),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd17)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[17]   )
    ,.unavailable_o       ( unavailable_o[17] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[17]   )
    ,.ipi_i               ( ipi_i[17]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[17*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile17_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile17_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_0_1_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_1_2_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_1_0_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_2_1_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_0_1_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_1_2_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_1_0_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_2_1_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_0_1_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_1_2_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_1_0_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_2_1_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_1_1_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_1_1_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_1_1_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_1_1_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_1_1_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_1_1_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_1_1_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_1_1_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_1_1_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_1_1_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_1_1_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_1_1_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_0_1_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_1_2_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_1_0_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_2_1_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_0_1_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_1_2_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_1_0_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_2_1_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_0_1_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_1_2_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_1_0_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_2_1_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_1_1_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_1_1_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_1_1_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_1_1_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_1_1_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_1_1_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_1_1_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_1_1_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_1_1_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_1_1_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_1_1_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_1_1_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_0_1_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_1_2_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_1_0_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_2_1_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_0_1_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_1_2_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_1_0_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_2_1_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_0_1_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_1_2_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_1_0_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_2_1_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_1_1_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_1_1_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_1_1_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_1_1_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_1_1_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_1_1_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_1_1_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_1_1_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_1_1_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_1_1_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_1_1_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_1_1_out_S_noc3_yummy )
);


tile
tile33 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[33] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd1),
    .default_coreid_y           (8'd2),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd33)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[33]   )
    ,.unavailable_o       ( unavailable_o[33] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[33]   )
    ,.ipi_i               ( ipi_i[33]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[33*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile33_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile33_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_1_1_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_2_2_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_2_0_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_3_1_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_1_1_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_2_2_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_2_0_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_3_1_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_1_1_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_2_2_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_2_0_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_3_1_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_2_1_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_2_1_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_2_1_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_2_1_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_2_1_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_2_1_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_2_1_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_2_1_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_2_1_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_2_1_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_2_1_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_2_1_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_1_1_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_2_2_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_2_0_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_3_1_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_1_1_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_2_2_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_2_0_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_3_1_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_1_1_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_2_2_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_2_0_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_3_1_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_2_1_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_2_1_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_2_1_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_2_1_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_2_1_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_2_1_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_2_1_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_2_1_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_2_1_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_2_1_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_2_1_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_2_1_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_1_1_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_2_2_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_2_0_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_3_1_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_1_1_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_2_2_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_2_0_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_3_1_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_1_1_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_2_2_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_2_0_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_3_1_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_2_1_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_2_1_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_2_1_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_2_1_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_2_1_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_2_1_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_2_1_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_2_1_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_2_1_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_2_1_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_2_1_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_2_1_out_S_noc3_yummy )
);


tile
tile49 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[49] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd1),
    .default_coreid_y           (8'd3),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd49)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[49]   )
    ,.unavailable_o       ( unavailable_o[49] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[49]   )
    ,.ipi_i               ( ipi_i[49]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[49*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile49_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile49_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_2_1_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_3_2_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_3_0_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_4_1_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_2_1_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_3_2_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_3_0_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_4_1_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_2_1_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_3_2_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_3_0_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_4_1_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_3_1_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_3_1_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_3_1_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_3_1_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_3_1_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_3_1_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_3_1_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_3_1_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_3_1_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_3_1_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_3_1_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_3_1_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_2_1_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_3_2_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_3_0_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_4_1_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_2_1_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_3_2_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_3_0_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_4_1_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_2_1_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_3_2_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_3_0_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_4_1_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_3_1_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_3_1_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_3_1_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_3_1_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_3_1_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_3_1_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_3_1_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_3_1_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_3_1_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_3_1_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_3_1_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_3_1_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_2_1_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_3_2_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_3_0_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_4_1_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_2_1_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_3_2_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_3_0_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_4_1_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_2_1_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_3_2_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_3_0_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_4_1_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_3_1_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_3_1_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_3_1_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_3_1_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_3_1_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_3_1_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_3_1_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_3_1_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_3_1_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_3_1_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_3_1_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_3_1_out_S_noc3_yummy )
);


tile
tile65 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[65] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd1),
    .default_coreid_y           (8'd4),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd65)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[65]   )
    ,.unavailable_o       ( unavailable_o[65] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[65]   )
    ,.ipi_i               ( ipi_i[65]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[65*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile65_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile65_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_3_1_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_4_2_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_4_0_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_5_1_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_3_1_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_4_2_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_4_0_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_5_1_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_3_1_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_4_2_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_4_0_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_5_1_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_4_1_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_4_1_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_4_1_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_4_1_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_4_1_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_4_1_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_4_1_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_4_1_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_4_1_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_4_1_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_4_1_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_4_1_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_3_1_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_4_2_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_4_0_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_5_1_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_3_1_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_4_2_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_4_0_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_5_1_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_3_1_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_4_2_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_4_0_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_5_1_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_4_1_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_4_1_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_4_1_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_4_1_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_4_1_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_4_1_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_4_1_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_4_1_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_4_1_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_4_1_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_4_1_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_4_1_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_3_1_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_4_2_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_4_0_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_5_1_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_3_1_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_4_2_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_4_0_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_5_1_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_3_1_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_4_2_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_4_0_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_5_1_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_4_1_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_4_1_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_4_1_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_4_1_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_4_1_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_4_1_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_4_1_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_4_1_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_4_1_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_4_1_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_4_1_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_4_1_out_S_noc3_yummy )
);


tile
tile81 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[81] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd1),
    .default_coreid_y           (8'd5),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd81)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[81]   )
    ,.unavailable_o       ( unavailable_o[81] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[81]   )
    ,.ipi_i               ( ipi_i[81]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[81*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile81_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile81_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_4_1_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_5_2_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_5_0_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_6_1_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_4_1_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_5_2_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_5_0_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_6_1_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_4_1_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_5_2_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_5_0_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_6_1_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_5_1_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_5_1_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_5_1_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_5_1_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_5_1_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_5_1_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_5_1_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_5_1_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_5_1_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_5_1_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_5_1_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_5_1_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_4_1_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_5_2_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_5_0_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_6_1_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_4_1_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_5_2_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_5_0_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_6_1_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_4_1_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_5_2_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_5_0_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_6_1_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_5_1_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_5_1_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_5_1_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_5_1_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_5_1_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_5_1_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_5_1_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_5_1_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_5_1_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_5_1_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_5_1_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_5_1_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_4_1_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_5_2_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_5_0_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_6_1_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_4_1_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_5_2_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_5_0_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_6_1_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_4_1_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_5_2_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_5_0_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_6_1_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_5_1_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_5_1_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_5_1_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_5_1_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_5_1_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_5_1_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_5_1_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_5_1_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_5_1_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_5_1_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_5_1_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_5_1_out_S_noc3_yummy )
);


tile
tile97 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[97] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd1),
    .default_coreid_y           (8'd6),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd97)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[97]   )
    ,.unavailable_o       ( unavailable_o[97] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[97]   )
    ,.ipi_i               ( ipi_i[97]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[97*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile97_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile97_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_5_1_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_6_2_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_6_0_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_7_1_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_5_1_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_6_2_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_6_0_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_7_1_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_5_1_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_6_2_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_6_0_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_7_1_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_6_1_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_6_1_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_6_1_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_6_1_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_6_1_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_6_1_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_6_1_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_6_1_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_6_1_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_6_1_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_6_1_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_6_1_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_5_1_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_6_2_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_6_0_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_7_1_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_5_1_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_6_2_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_6_0_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_7_1_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_5_1_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_6_2_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_6_0_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_7_1_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_6_1_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_6_1_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_6_1_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_6_1_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_6_1_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_6_1_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_6_1_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_6_1_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_6_1_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_6_1_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_6_1_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_6_1_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_5_1_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_6_2_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_6_0_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_7_1_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_5_1_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_6_2_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_6_0_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_7_1_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_5_1_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_6_2_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_6_0_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_7_1_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_6_1_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_6_1_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_6_1_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_6_1_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_6_1_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_6_1_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_6_1_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_6_1_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_6_1_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_6_1_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_6_1_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_6_1_out_S_noc3_yummy )
);


tile
tile113 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[113] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd1),
    .default_coreid_y           (8'd7),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd113)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[113]   )
    ,.unavailable_o       ( unavailable_o[113] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[113]   )
    ,.ipi_i               ( ipi_i[113]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[113*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile113_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile113_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_6_1_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_7_2_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_7_0_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_8_1_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_6_1_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_7_2_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_7_0_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_8_1_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_6_1_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_7_2_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_7_0_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_8_1_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_7_1_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_7_1_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_7_1_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_7_1_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_7_1_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_7_1_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_7_1_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_7_1_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_7_1_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_7_1_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_7_1_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_7_1_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_6_1_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_7_2_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_7_0_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_8_1_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_6_1_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_7_2_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_7_0_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_8_1_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_6_1_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_7_2_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_7_0_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_8_1_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_7_1_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_7_1_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_7_1_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_7_1_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_7_1_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_7_1_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_7_1_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_7_1_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_7_1_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_7_1_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_7_1_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_7_1_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_6_1_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_7_2_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_7_0_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_8_1_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_6_1_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_7_2_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_7_0_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_8_1_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_6_1_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_7_2_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_7_0_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_8_1_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_7_1_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_7_1_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_7_1_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_7_1_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_7_1_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_7_1_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_7_1_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_7_1_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_7_1_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_7_1_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_7_1_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_7_1_out_S_noc3_yummy )
);


tile
tile129 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[129] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd1),
    .default_coreid_y           (8'd8),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd129)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[129]   )
    ,.unavailable_o       ( unavailable_o[129] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[129]   )
    ,.ipi_i               ( ipi_i[129]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[129*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile129_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile129_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_7_1_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_8_2_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_8_0_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_9_1_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_7_1_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_8_2_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_8_0_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_9_1_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_7_1_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_8_2_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_8_0_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_9_1_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_8_1_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_8_1_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_8_1_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_8_1_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_8_1_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_8_1_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_8_1_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_8_1_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_8_1_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_8_1_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_8_1_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_8_1_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_7_1_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_8_2_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_8_0_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_9_1_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_7_1_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_8_2_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_8_0_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_9_1_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_7_1_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_8_2_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_8_0_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_9_1_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_8_1_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_8_1_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_8_1_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_8_1_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_8_1_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_8_1_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_8_1_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_8_1_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_8_1_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_8_1_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_8_1_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_8_1_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_7_1_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_8_2_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_8_0_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_9_1_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_7_1_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_8_2_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_8_0_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_9_1_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_7_1_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_8_2_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_8_0_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_9_1_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_8_1_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_8_1_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_8_1_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_8_1_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_8_1_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_8_1_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_8_1_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_8_1_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_8_1_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_8_1_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_8_1_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_8_1_out_S_noc3_yummy )
);


tile
tile145 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[145] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd1),
    .default_coreid_y           (8'd9),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd145)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[145]   )
    ,.unavailable_o       ( unavailable_o[145] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[145]   )
    ,.ipi_i               ( ipi_i[145]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[145*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile145_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile145_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_8_1_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_9_2_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_9_0_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_10_1_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_8_1_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_9_2_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_9_0_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_10_1_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_8_1_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_9_2_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_9_0_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_10_1_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_9_1_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_9_1_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_9_1_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_9_1_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_9_1_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_9_1_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_9_1_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_9_1_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_9_1_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_9_1_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_9_1_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_9_1_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_8_1_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_9_2_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_9_0_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_10_1_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_8_1_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_9_2_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_9_0_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_10_1_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_8_1_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_9_2_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_9_0_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_10_1_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_9_1_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_9_1_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_9_1_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_9_1_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_9_1_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_9_1_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_9_1_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_9_1_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_9_1_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_9_1_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_9_1_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_9_1_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_8_1_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_9_2_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_9_0_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_10_1_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_8_1_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_9_2_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_9_0_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_10_1_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_8_1_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_9_2_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_9_0_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_10_1_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_9_1_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_9_1_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_9_1_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_9_1_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_9_1_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_9_1_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_9_1_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_9_1_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_9_1_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_9_1_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_9_1_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_9_1_out_S_noc3_yummy )
);


tile
tile161 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[161] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd1),
    .default_coreid_y           (8'd10),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd161)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[161]   )
    ,.unavailable_o       ( unavailable_o[161] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[161]   )
    ,.ipi_i               ( ipi_i[161]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[161*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile161_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile161_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_9_1_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_10_2_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_10_0_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_11_1_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_9_1_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_10_2_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_10_0_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_11_1_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_9_1_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_10_2_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_10_0_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_11_1_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_10_1_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_10_1_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_10_1_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_10_1_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_10_1_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_10_1_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_10_1_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_10_1_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_10_1_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_10_1_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_10_1_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_10_1_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_9_1_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_10_2_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_10_0_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_11_1_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_9_1_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_10_2_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_10_0_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_11_1_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_9_1_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_10_2_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_10_0_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_11_1_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_10_1_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_10_1_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_10_1_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_10_1_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_10_1_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_10_1_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_10_1_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_10_1_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_10_1_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_10_1_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_10_1_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_10_1_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_9_1_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_10_2_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_10_0_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_11_1_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_9_1_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_10_2_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_10_0_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_11_1_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_9_1_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_10_2_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_10_0_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_11_1_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_10_1_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_10_1_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_10_1_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_10_1_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_10_1_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_10_1_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_10_1_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_10_1_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_10_1_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_10_1_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_10_1_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_10_1_out_S_noc3_yummy )
);


tile
tile177 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[177] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd1),
    .default_coreid_y           (8'd11),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd177)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[177]   )
    ,.unavailable_o       ( unavailable_o[177] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[177]   )
    ,.ipi_i               ( ipi_i[177]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[177*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile177_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile177_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_10_1_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_11_2_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_11_0_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_12_1_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_10_1_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_11_2_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_11_0_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_12_1_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_10_1_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_11_2_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_11_0_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_12_1_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_11_1_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_11_1_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_11_1_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_11_1_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_11_1_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_11_1_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_11_1_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_11_1_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_11_1_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_11_1_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_11_1_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_11_1_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_10_1_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_11_2_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_11_0_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_12_1_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_10_1_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_11_2_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_11_0_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_12_1_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_10_1_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_11_2_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_11_0_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_12_1_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_11_1_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_11_1_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_11_1_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_11_1_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_11_1_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_11_1_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_11_1_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_11_1_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_11_1_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_11_1_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_11_1_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_11_1_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_10_1_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_11_2_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_11_0_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_12_1_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_10_1_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_11_2_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_11_0_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_12_1_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_10_1_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_11_2_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_11_0_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_12_1_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_11_1_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_11_1_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_11_1_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_11_1_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_11_1_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_11_1_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_11_1_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_11_1_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_11_1_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_11_1_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_11_1_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_11_1_out_S_noc3_yummy )
);


tile
tile193 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[193] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd1),
    .default_coreid_y           (8'd12),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd193)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[193]   )
    ,.unavailable_o       ( unavailable_o[193] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[193]   )
    ,.ipi_i               ( ipi_i[193]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[193*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile193_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile193_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_11_1_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_12_2_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_12_0_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_13_1_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_11_1_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_12_2_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_12_0_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_13_1_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_11_1_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_12_2_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_12_0_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_13_1_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_12_1_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_12_1_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_12_1_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_12_1_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_12_1_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_12_1_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_12_1_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_12_1_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_12_1_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_12_1_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_12_1_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_12_1_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_11_1_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_12_2_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_12_0_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_13_1_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_11_1_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_12_2_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_12_0_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_13_1_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_11_1_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_12_2_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_12_0_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_13_1_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_12_1_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_12_1_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_12_1_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_12_1_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_12_1_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_12_1_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_12_1_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_12_1_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_12_1_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_12_1_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_12_1_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_12_1_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_11_1_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_12_2_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_12_0_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_13_1_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_11_1_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_12_2_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_12_0_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_13_1_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_11_1_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_12_2_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_12_0_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_13_1_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_12_1_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_12_1_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_12_1_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_12_1_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_12_1_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_12_1_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_12_1_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_12_1_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_12_1_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_12_1_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_12_1_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_12_1_out_S_noc3_yummy )
);


tile
tile209 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[209] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd1),
    .default_coreid_y           (8'd13),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd209)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[209]   )
    ,.unavailable_o       ( unavailable_o[209] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[209]   )
    ,.ipi_i               ( ipi_i[209]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[209*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile209_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile209_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_12_1_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_13_2_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_13_0_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_14_1_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_12_1_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_13_2_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_13_0_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_14_1_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_12_1_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_13_2_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_13_0_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_14_1_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_13_1_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_13_1_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_13_1_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_13_1_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_13_1_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_13_1_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_13_1_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_13_1_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_13_1_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_13_1_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_13_1_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_13_1_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_12_1_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_13_2_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_13_0_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_14_1_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_12_1_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_13_2_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_13_0_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_14_1_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_12_1_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_13_2_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_13_0_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_14_1_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_13_1_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_13_1_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_13_1_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_13_1_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_13_1_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_13_1_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_13_1_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_13_1_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_13_1_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_13_1_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_13_1_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_13_1_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_12_1_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_13_2_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_13_0_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_14_1_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_12_1_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_13_2_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_13_0_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_14_1_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_12_1_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_13_2_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_13_0_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_14_1_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_13_1_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_13_1_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_13_1_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_13_1_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_13_1_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_13_1_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_13_1_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_13_1_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_13_1_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_13_1_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_13_1_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_13_1_out_S_noc3_yummy )
);


tile
tile225 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[225] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd1),
    .default_coreid_y           (8'd14),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd225)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[225]   )
    ,.unavailable_o       ( unavailable_o[225] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[225]   )
    ,.ipi_i               ( ipi_i[225]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[225*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile225_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile225_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_13_1_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_14_2_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_14_0_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_15_1_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_13_1_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_14_2_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_14_0_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_15_1_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_13_1_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_14_2_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_14_0_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_15_1_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_14_1_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_14_1_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_14_1_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_14_1_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_14_1_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_14_1_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_14_1_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_14_1_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_14_1_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_14_1_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_14_1_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_14_1_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_13_1_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_14_2_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_14_0_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_15_1_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_13_1_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_14_2_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_14_0_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_15_1_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_13_1_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_14_2_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_14_0_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_15_1_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_14_1_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_14_1_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_14_1_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_14_1_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_14_1_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_14_1_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_14_1_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_14_1_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_14_1_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_14_1_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_14_1_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_14_1_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_13_1_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_14_2_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_14_0_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_15_1_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_13_1_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_14_2_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_14_0_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_15_1_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_13_1_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_14_2_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_14_0_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_15_1_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_14_1_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_14_1_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_14_1_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_14_1_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_14_1_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_14_1_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_14_1_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_14_1_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_14_1_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_14_1_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_14_1_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_14_1_out_S_noc3_yummy )
);


tile
tile241 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[241] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd1),
    .default_coreid_y           (8'd15),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd241)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[241]   )
    ,.unavailable_o       ( unavailable_o[241] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[241]   )
    ,.ipi_i               ( ipi_i[241]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[241*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile241_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile241_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_14_1_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_15_2_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_15_0_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( dummy_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_14_1_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_15_2_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_15_0_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( dummy_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_14_1_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_15_2_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_15_0_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( dummy_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_15_1_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_15_1_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_15_1_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_15_1_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_15_1_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_15_1_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_15_1_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_15_1_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_15_1_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_15_1_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_15_1_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_15_1_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_14_1_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_15_2_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_15_0_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( dummy_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_14_1_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_15_2_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_15_0_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( dummy_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_14_1_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_15_2_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_15_0_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( dummy_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_15_1_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_15_1_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_15_1_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_15_1_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_15_1_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_15_1_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_15_1_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_15_1_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_15_1_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_15_1_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_15_1_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_15_1_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_14_1_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_15_2_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_15_0_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( dummy_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_14_1_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_15_2_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_15_0_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( dummy_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_14_1_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_15_2_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_15_0_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( dummy_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_15_1_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_15_1_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_15_1_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_15_1_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_15_1_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_15_1_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_15_1_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_15_1_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_15_1_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_15_1_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_15_1_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_15_1_out_S_noc3_yummy )
);


tile
tile2 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[2] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd2),
    .default_coreid_y           (8'd0),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd2)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[2]   )
    ,.unavailable_o       ( unavailable_o[2] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[2]   )
    ,.ipi_i               ( ipi_i[2]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[2*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile2_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile2_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( dummy_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_0_3_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_0_1_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_1_2_out_N_noc1_data   ),
    .dyn0_validIn_N      ( dummy_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_0_3_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_0_1_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_1_2_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( dummy_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_0_3_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_0_1_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_1_2_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_0_2_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_0_2_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_0_2_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_0_2_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_0_2_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_0_2_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_0_2_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_0_2_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_0_2_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_0_2_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_0_2_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_0_2_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( dummy_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_0_3_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_0_1_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_1_2_out_N_noc2_data   ),
    .dyn1_validIn_N      ( dummy_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_0_3_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_0_1_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_1_2_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( dummy_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_0_3_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_0_1_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_1_2_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_0_2_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_0_2_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_0_2_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_0_2_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_0_2_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_0_2_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_0_2_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_0_2_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_0_2_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_0_2_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_0_2_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_0_2_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( dummy_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_0_3_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_0_1_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_1_2_out_N_noc3_data   ),
    .dyn2_validIn_N      ( dummy_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_0_3_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_0_1_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_1_2_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( dummy_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_0_3_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_0_1_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_1_2_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_0_2_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_0_2_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_0_2_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_0_2_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_0_2_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_0_2_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_0_2_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_0_2_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_0_2_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_0_2_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_0_2_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_0_2_out_S_noc3_yummy )
);


tile
tile18 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[18] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd2),
    .default_coreid_y           (8'd1),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd18)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[18]   )
    ,.unavailable_o       ( unavailable_o[18] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[18]   )
    ,.ipi_i               ( ipi_i[18]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[18*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile18_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile18_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_0_2_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_1_3_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_1_1_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_2_2_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_0_2_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_1_3_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_1_1_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_2_2_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_0_2_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_1_3_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_1_1_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_2_2_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_1_2_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_1_2_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_1_2_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_1_2_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_1_2_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_1_2_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_1_2_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_1_2_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_1_2_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_1_2_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_1_2_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_1_2_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_0_2_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_1_3_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_1_1_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_2_2_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_0_2_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_1_3_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_1_1_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_2_2_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_0_2_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_1_3_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_1_1_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_2_2_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_1_2_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_1_2_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_1_2_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_1_2_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_1_2_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_1_2_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_1_2_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_1_2_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_1_2_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_1_2_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_1_2_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_1_2_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_0_2_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_1_3_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_1_1_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_2_2_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_0_2_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_1_3_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_1_1_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_2_2_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_0_2_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_1_3_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_1_1_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_2_2_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_1_2_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_1_2_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_1_2_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_1_2_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_1_2_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_1_2_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_1_2_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_1_2_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_1_2_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_1_2_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_1_2_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_1_2_out_S_noc3_yummy )
);


tile
tile34 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[34] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd2),
    .default_coreid_y           (8'd2),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd34)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[34]   )
    ,.unavailable_o       ( unavailable_o[34] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[34]   )
    ,.ipi_i               ( ipi_i[34]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[34*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile34_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile34_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_1_2_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_2_3_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_2_1_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_3_2_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_1_2_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_2_3_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_2_1_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_3_2_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_1_2_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_2_3_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_2_1_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_3_2_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_2_2_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_2_2_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_2_2_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_2_2_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_2_2_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_2_2_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_2_2_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_2_2_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_2_2_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_2_2_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_2_2_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_2_2_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_1_2_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_2_3_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_2_1_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_3_2_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_1_2_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_2_3_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_2_1_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_3_2_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_1_2_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_2_3_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_2_1_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_3_2_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_2_2_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_2_2_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_2_2_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_2_2_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_2_2_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_2_2_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_2_2_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_2_2_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_2_2_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_2_2_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_2_2_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_2_2_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_1_2_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_2_3_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_2_1_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_3_2_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_1_2_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_2_3_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_2_1_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_3_2_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_1_2_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_2_3_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_2_1_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_3_2_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_2_2_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_2_2_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_2_2_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_2_2_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_2_2_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_2_2_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_2_2_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_2_2_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_2_2_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_2_2_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_2_2_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_2_2_out_S_noc3_yummy )
);


tile
tile50 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[50] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd2),
    .default_coreid_y           (8'd3),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd50)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[50]   )
    ,.unavailable_o       ( unavailable_o[50] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[50]   )
    ,.ipi_i               ( ipi_i[50]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[50*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile50_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile50_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_2_2_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_3_3_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_3_1_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_4_2_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_2_2_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_3_3_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_3_1_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_4_2_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_2_2_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_3_3_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_3_1_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_4_2_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_3_2_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_3_2_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_3_2_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_3_2_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_3_2_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_3_2_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_3_2_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_3_2_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_3_2_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_3_2_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_3_2_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_3_2_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_2_2_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_3_3_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_3_1_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_4_2_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_2_2_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_3_3_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_3_1_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_4_2_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_2_2_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_3_3_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_3_1_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_4_2_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_3_2_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_3_2_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_3_2_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_3_2_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_3_2_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_3_2_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_3_2_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_3_2_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_3_2_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_3_2_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_3_2_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_3_2_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_2_2_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_3_3_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_3_1_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_4_2_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_2_2_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_3_3_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_3_1_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_4_2_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_2_2_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_3_3_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_3_1_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_4_2_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_3_2_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_3_2_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_3_2_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_3_2_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_3_2_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_3_2_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_3_2_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_3_2_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_3_2_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_3_2_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_3_2_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_3_2_out_S_noc3_yummy )
);


tile
tile66 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[66] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd2),
    .default_coreid_y           (8'd4),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd66)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[66]   )
    ,.unavailable_o       ( unavailable_o[66] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[66]   )
    ,.ipi_i               ( ipi_i[66]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[66*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile66_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile66_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_3_2_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_4_3_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_4_1_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_5_2_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_3_2_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_4_3_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_4_1_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_5_2_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_3_2_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_4_3_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_4_1_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_5_2_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_4_2_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_4_2_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_4_2_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_4_2_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_4_2_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_4_2_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_4_2_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_4_2_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_4_2_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_4_2_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_4_2_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_4_2_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_3_2_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_4_3_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_4_1_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_5_2_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_3_2_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_4_3_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_4_1_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_5_2_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_3_2_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_4_3_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_4_1_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_5_2_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_4_2_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_4_2_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_4_2_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_4_2_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_4_2_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_4_2_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_4_2_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_4_2_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_4_2_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_4_2_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_4_2_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_4_2_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_3_2_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_4_3_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_4_1_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_5_2_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_3_2_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_4_3_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_4_1_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_5_2_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_3_2_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_4_3_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_4_1_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_5_2_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_4_2_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_4_2_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_4_2_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_4_2_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_4_2_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_4_2_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_4_2_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_4_2_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_4_2_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_4_2_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_4_2_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_4_2_out_S_noc3_yummy )
);


tile
tile82 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[82] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd2),
    .default_coreid_y           (8'd5),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd82)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[82]   )
    ,.unavailable_o       ( unavailable_o[82] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[82]   )
    ,.ipi_i               ( ipi_i[82]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[82*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile82_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile82_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_4_2_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_5_3_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_5_1_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_6_2_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_4_2_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_5_3_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_5_1_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_6_2_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_4_2_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_5_3_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_5_1_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_6_2_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_5_2_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_5_2_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_5_2_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_5_2_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_5_2_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_5_2_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_5_2_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_5_2_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_5_2_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_5_2_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_5_2_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_5_2_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_4_2_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_5_3_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_5_1_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_6_2_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_4_2_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_5_3_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_5_1_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_6_2_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_4_2_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_5_3_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_5_1_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_6_2_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_5_2_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_5_2_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_5_2_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_5_2_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_5_2_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_5_2_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_5_2_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_5_2_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_5_2_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_5_2_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_5_2_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_5_2_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_4_2_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_5_3_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_5_1_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_6_2_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_4_2_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_5_3_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_5_1_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_6_2_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_4_2_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_5_3_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_5_1_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_6_2_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_5_2_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_5_2_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_5_2_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_5_2_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_5_2_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_5_2_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_5_2_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_5_2_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_5_2_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_5_2_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_5_2_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_5_2_out_S_noc3_yummy )
);


tile
tile98 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[98] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd2),
    .default_coreid_y           (8'd6),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd98)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[98]   )
    ,.unavailable_o       ( unavailable_o[98] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[98]   )
    ,.ipi_i               ( ipi_i[98]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[98*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile98_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile98_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_5_2_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_6_3_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_6_1_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_7_2_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_5_2_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_6_3_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_6_1_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_7_2_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_5_2_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_6_3_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_6_1_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_7_2_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_6_2_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_6_2_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_6_2_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_6_2_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_6_2_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_6_2_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_6_2_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_6_2_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_6_2_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_6_2_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_6_2_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_6_2_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_5_2_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_6_3_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_6_1_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_7_2_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_5_2_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_6_3_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_6_1_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_7_2_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_5_2_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_6_3_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_6_1_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_7_2_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_6_2_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_6_2_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_6_2_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_6_2_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_6_2_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_6_2_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_6_2_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_6_2_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_6_2_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_6_2_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_6_2_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_6_2_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_5_2_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_6_3_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_6_1_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_7_2_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_5_2_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_6_3_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_6_1_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_7_2_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_5_2_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_6_3_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_6_1_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_7_2_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_6_2_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_6_2_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_6_2_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_6_2_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_6_2_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_6_2_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_6_2_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_6_2_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_6_2_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_6_2_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_6_2_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_6_2_out_S_noc3_yummy )
);


tile
tile114 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[114] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd2),
    .default_coreid_y           (8'd7),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd114)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[114]   )
    ,.unavailable_o       ( unavailable_o[114] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[114]   )
    ,.ipi_i               ( ipi_i[114]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[114*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile114_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile114_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_6_2_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_7_3_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_7_1_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_8_2_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_6_2_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_7_3_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_7_1_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_8_2_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_6_2_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_7_3_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_7_1_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_8_2_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_7_2_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_7_2_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_7_2_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_7_2_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_7_2_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_7_2_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_7_2_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_7_2_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_7_2_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_7_2_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_7_2_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_7_2_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_6_2_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_7_3_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_7_1_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_8_2_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_6_2_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_7_3_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_7_1_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_8_2_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_6_2_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_7_3_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_7_1_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_8_2_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_7_2_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_7_2_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_7_2_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_7_2_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_7_2_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_7_2_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_7_2_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_7_2_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_7_2_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_7_2_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_7_2_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_7_2_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_6_2_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_7_3_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_7_1_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_8_2_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_6_2_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_7_3_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_7_1_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_8_2_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_6_2_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_7_3_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_7_1_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_8_2_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_7_2_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_7_2_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_7_2_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_7_2_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_7_2_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_7_2_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_7_2_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_7_2_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_7_2_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_7_2_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_7_2_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_7_2_out_S_noc3_yummy )
);


tile
tile130 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[130] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd2),
    .default_coreid_y           (8'd8),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd130)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[130]   )
    ,.unavailable_o       ( unavailable_o[130] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[130]   )
    ,.ipi_i               ( ipi_i[130]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[130*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile130_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile130_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_7_2_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_8_3_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_8_1_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_9_2_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_7_2_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_8_3_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_8_1_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_9_2_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_7_2_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_8_3_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_8_1_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_9_2_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_8_2_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_8_2_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_8_2_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_8_2_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_8_2_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_8_2_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_8_2_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_8_2_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_8_2_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_8_2_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_8_2_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_8_2_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_7_2_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_8_3_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_8_1_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_9_2_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_7_2_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_8_3_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_8_1_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_9_2_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_7_2_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_8_3_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_8_1_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_9_2_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_8_2_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_8_2_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_8_2_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_8_2_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_8_2_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_8_2_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_8_2_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_8_2_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_8_2_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_8_2_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_8_2_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_8_2_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_7_2_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_8_3_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_8_1_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_9_2_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_7_2_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_8_3_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_8_1_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_9_2_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_7_2_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_8_3_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_8_1_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_9_2_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_8_2_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_8_2_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_8_2_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_8_2_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_8_2_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_8_2_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_8_2_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_8_2_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_8_2_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_8_2_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_8_2_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_8_2_out_S_noc3_yummy )
);


tile
tile146 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[146] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd2),
    .default_coreid_y           (8'd9),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd146)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[146]   )
    ,.unavailable_o       ( unavailable_o[146] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[146]   )
    ,.ipi_i               ( ipi_i[146]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[146*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile146_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile146_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_8_2_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_9_3_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_9_1_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_10_2_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_8_2_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_9_3_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_9_1_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_10_2_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_8_2_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_9_3_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_9_1_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_10_2_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_9_2_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_9_2_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_9_2_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_9_2_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_9_2_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_9_2_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_9_2_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_9_2_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_9_2_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_9_2_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_9_2_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_9_2_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_8_2_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_9_3_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_9_1_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_10_2_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_8_2_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_9_3_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_9_1_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_10_2_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_8_2_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_9_3_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_9_1_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_10_2_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_9_2_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_9_2_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_9_2_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_9_2_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_9_2_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_9_2_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_9_2_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_9_2_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_9_2_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_9_2_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_9_2_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_9_2_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_8_2_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_9_3_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_9_1_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_10_2_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_8_2_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_9_3_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_9_1_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_10_2_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_8_2_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_9_3_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_9_1_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_10_2_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_9_2_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_9_2_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_9_2_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_9_2_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_9_2_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_9_2_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_9_2_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_9_2_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_9_2_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_9_2_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_9_2_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_9_2_out_S_noc3_yummy )
);


tile
tile162 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[162] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd2),
    .default_coreid_y           (8'd10),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd162)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[162]   )
    ,.unavailable_o       ( unavailable_o[162] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[162]   )
    ,.ipi_i               ( ipi_i[162]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[162*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile162_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile162_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_9_2_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_10_3_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_10_1_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_11_2_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_9_2_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_10_3_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_10_1_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_11_2_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_9_2_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_10_3_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_10_1_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_11_2_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_10_2_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_10_2_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_10_2_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_10_2_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_10_2_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_10_2_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_10_2_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_10_2_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_10_2_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_10_2_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_10_2_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_10_2_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_9_2_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_10_3_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_10_1_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_11_2_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_9_2_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_10_3_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_10_1_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_11_2_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_9_2_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_10_3_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_10_1_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_11_2_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_10_2_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_10_2_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_10_2_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_10_2_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_10_2_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_10_2_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_10_2_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_10_2_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_10_2_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_10_2_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_10_2_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_10_2_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_9_2_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_10_3_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_10_1_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_11_2_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_9_2_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_10_3_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_10_1_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_11_2_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_9_2_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_10_3_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_10_1_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_11_2_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_10_2_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_10_2_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_10_2_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_10_2_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_10_2_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_10_2_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_10_2_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_10_2_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_10_2_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_10_2_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_10_2_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_10_2_out_S_noc3_yummy )
);


tile
tile178 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[178] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd2),
    .default_coreid_y           (8'd11),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd178)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[178]   )
    ,.unavailable_o       ( unavailable_o[178] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[178]   )
    ,.ipi_i               ( ipi_i[178]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[178*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile178_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile178_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_10_2_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_11_3_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_11_1_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_12_2_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_10_2_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_11_3_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_11_1_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_12_2_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_10_2_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_11_3_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_11_1_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_12_2_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_11_2_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_11_2_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_11_2_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_11_2_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_11_2_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_11_2_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_11_2_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_11_2_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_11_2_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_11_2_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_11_2_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_11_2_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_10_2_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_11_3_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_11_1_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_12_2_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_10_2_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_11_3_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_11_1_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_12_2_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_10_2_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_11_3_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_11_1_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_12_2_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_11_2_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_11_2_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_11_2_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_11_2_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_11_2_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_11_2_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_11_2_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_11_2_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_11_2_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_11_2_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_11_2_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_11_2_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_10_2_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_11_3_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_11_1_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_12_2_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_10_2_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_11_3_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_11_1_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_12_2_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_10_2_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_11_3_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_11_1_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_12_2_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_11_2_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_11_2_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_11_2_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_11_2_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_11_2_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_11_2_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_11_2_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_11_2_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_11_2_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_11_2_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_11_2_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_11_2_out_S_noc3_yummy )
);


tile
tile194 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[194] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd2),
    .default_coreid_y           (8'd12),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd194)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[194]   )
    ,.unavailable_o       ( unavailable_o[194] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[194]   )
    ,.ipi_i               ( ipi_i[194]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[194*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile194_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile194_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_11_2_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_12_3_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_12_1_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_13_2_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_11_2_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_12_3_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_12_1_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_13_2_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_11_2_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_12_3_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_12_1_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_13_2_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_12_2_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_12_2_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_12_2_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_12_2_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_12_2_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_12_2_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_12_2_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_12_2_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_12_2_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_12_2_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_12_2_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_12_2_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_11_2_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_12_3_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_12_1_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_13_2_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_11_2_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_12_3_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_12_1_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_13_2_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_11_2_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_12_3_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_12_1_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_13_2_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_12_2_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_12_2_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_12_2_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_12_2_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_12_2_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_12_2_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_12_2_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_12_2_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_12_2_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_12_2_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_12_2_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_12_2_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_11_2_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_12_3_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_12_1_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_13_2_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_11_2_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_12_3_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_12_1_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_13_2_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_11_2_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_12_3_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_12_1_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_13_2_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_12_2_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_12_2_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_12_2_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_12_2_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_12_2_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_12_2_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_12_2_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_12_2_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_12_2_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_12_2_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_12_2_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_12_2_out_S_noc3_yummy )
);


tile
tile210 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[210] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd2),
    .default_coreid_y           (8'd13),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd210)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[210]   )
    ,.unavailable_o       ( unavailable_o[210] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[210]   )
    ,.ipi_i               ( ipi_i[210]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[210*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile210_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile210_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_12_2_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_13_3_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_13_1_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_14_2_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_12_2_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_13_3_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_13_1_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_14_2_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_12_2_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_13_3_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_13_1_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_14_2_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_13_2_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_13_2_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_13_2_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_13_2_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_13_2_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_13_2_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_13_2_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_13_2_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_13_2_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_13_2_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_13_2_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_13_2_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_12_2_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_13_3_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_13_1_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_14_2_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_12_2_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_13_3_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_13_1_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_14_2_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_12_2_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_13_3_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_13_1_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_14_2_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_13_2_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_13_2_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_13_2_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_13_2_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_13_2_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_13_2_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_13_2_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_13_2_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_13_2_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_13_2_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_13_2_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_13_2_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_12_2_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_13_3_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_13_1_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_14_2_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_12_2_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_13_3_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_13_1_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_14_2_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_12_2_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_13_3_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_13_1_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_14_2_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_13_2_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_13_2_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_13_2_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_13_2_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_13_2_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_13_2_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_13_2_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_13_2_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_13_2_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_13_2_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_13_2_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_13_2_out_S_noc3_yummy )
);


tile
tile226 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[226] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd2),
    .default_coreid_y           (8'd14),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd226)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[226]   )
    ,.unavailable_o       ( unavailable_o[226] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[226]   )
    ,.ipi_i               ( ipi_i[226]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[226*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile226_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile226_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_13_2_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_14_3_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_14_1_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_15_2_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_13_2_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_14_3_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_14_1_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_15_2_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_13_2_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_14_3_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_14_1_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_15_2_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_14_2_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_14_2_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_14_2_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_14_2_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_14_2_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_14_2_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_14_2_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_14_2_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_14_2_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_14_2_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_14_2_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_14_2_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_13_2_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_14_3_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_14_1_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_15_2_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_13_2_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_14_3_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_14_1_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_15_2_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_13_2_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_14_3_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_14_1_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_15_2_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_14_2_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_14_2_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_14_2_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_14_2_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_14_2_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_14_2_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_14_2_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_14_2_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_14_2_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_14_2_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_14_2_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_14_2_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_13_2_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_14_3_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_14_1_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_15_2_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_13_2_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_14_3_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_14_1_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_15_2_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_13_2_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_14_3_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_14_1_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_15_2_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_14_2_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_14_2_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_14_2_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_14_2_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_14_2_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_14_2_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_14_2_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_14_2_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_14_2_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_14_2_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_14_2_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_14_2_out_S_noc3_yummy )
);


tile
tile242 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[242] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd2),
    .default_coreid_y           (8'd15),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd242)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[242]   )
    ,.unavailable_o       ( unavailable_o[242] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[242]   )
    ,.ipi_i               ( ipi_i[242]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[242*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile242_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile242_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_14_2_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_15_3_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_15_1_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( dummy_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_14_2_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_15_3_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_15_1_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( dummy_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_14_2_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_15_3_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_15_1_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( dummy_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_15_2_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_15_2_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_15_2_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_15_2_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_15_2_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_15_2_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_15_2_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_15_2_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_15_2_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_15_2_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_15_2_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_15_2_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_14_2_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_15_3_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_15_1_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( dummy_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_14_2_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_15_3_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_15_1_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( dummy_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_14_2_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_15_3_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_15_1_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( dummy_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_15_2_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_15_2_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_15_2_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_15_2_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_15_2_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_15_2_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_15_2_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_15_2_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_15_2_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_15_2_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_15_2_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_15_2_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_14_2_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_15_3_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_15_1_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( dummy_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_14_2_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_15_3_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_15_1_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( dummy_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_14_2_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_15_3_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_15_1_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( dummy_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_15_2_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_15_2_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_15_2_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_15_2_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_15_2_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_15_2_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_15_2_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_15_2_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_15_2_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_15_2_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_15_2_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_15_2_out_S_noc3_yummy )
);


tile
tile3 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[3] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd3),
    .default_coreid_y           (8'd0),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd3)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[3]   )
    ,.unavailable_o       ( unavailable_o[3] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[3]   )
    ,.ipi_i               ( ipi_i[3]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[3*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile3_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile3_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( dummy_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_0_4_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_0_2_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_1_3_out_N_noc1_data   ),
    .dyn0_validIn_N      ( dummy_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_0_4_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_0_2_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_1_3_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( dummy_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_0_4_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_0_2_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_1_3_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_0_3_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_0_3_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_0_3_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_0_3_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_0_3_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_0_3_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_0_3_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_0_3_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_0_3_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_0_3_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_0_3_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_0_3_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( dummy_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_0_4_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_0_2_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_1_3_out_N_noc2_data   ),
    .dyn1_validIn_N      ( dummy_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_0_4_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_0_2_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_1_3_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( dummy_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_0_4_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_0_2_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_1_3_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_0_3_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_0_3_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_0_3_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_0_3_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_0_3_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_0_3_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_0_3_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_0_3_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_0_3_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_0_3_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_0_3_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_0_3_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( dummy_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_0_4_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_0_2_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_1_3_out_N_noc3_data   ),
    .dyn2_validIn_N      ( dummy_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_0_4_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_0_2_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_1_3_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( dummy_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_0_4_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_0_2_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_1_3_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_0_3_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_0_3_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_0_3_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_0_3_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_0_3_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_0_3_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_0_3_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_0_3_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_0_3_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_0_3_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_0_3_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_0_3_out_S_noc3_yummy )
);


tile
tile19 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[19] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd3),
    .default_coreid_y           (8'd1),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd19)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[19]   )
    ,.unavailable_o       ( unavailable_o[19] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[19]   )
    ,.ipi_i               ( ipi_i[19]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[19*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile19_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile19_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_0_3_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_1_4_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_1_2_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_2_3_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_0_3_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_1_4_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_1_2_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_2_3_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_0_3_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_1_4_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_1_2_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_2_3_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_1_3_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_1_3_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_1_3_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_1_3_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_1_3_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_1_3_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_1_3_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_1_3_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_1_3_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_1_3_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_1_3_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_1_3_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_0_3_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_1_4_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_1_2_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_2_3_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_0_3_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_1_4_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_1_2_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_2_3_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_0_3_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_1_4_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_1_2_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_2_3_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_1_3_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_1_3_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_1_3_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_1_3_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_1_3_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_1_3_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_1_3_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_1_3_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_1_3_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_1_3_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_1_3_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_1_3_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_0_3_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_1_4_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_1_2_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_2_3_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_0_3_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_1_4_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_1_2_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_2_3_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_0_3_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_1_4_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_1_2_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_2_3_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_1_3_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_1_3_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_1_3_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_1_3_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_1_3_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_1_3_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_1_3_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_1_3_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_1_3_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_1_3_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_1_3_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_1_3_out_S_noc3_yummy )
);


tile
tile35 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[35] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd3),
    .default_coreid_y           (8'd2),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd35)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[35]   )
    ,.unavailable_o       ( unavailable_o[35] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[35]   )
    ,.ipi_i               ( ipi_i[35]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[35*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile35_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile35_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_1_3_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_2_4_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_2_2_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_3_3_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_1_3_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_2_4_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_2_2_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_3_3_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_1_3_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_2_4_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_2_2_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_3_3_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_2_3_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_2_3_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_2_3_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_2_3_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_2_3_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_2_3_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_2_3_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_2_3_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_2_3_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_2_3_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_2_3_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_2_3_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_1_3_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_2_4_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_2_2_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_3_3_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_1_3_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_2_4_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_2_2_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_3_3_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_1_3_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_2_4_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_2_2_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_3_3_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_2_3_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_2_3_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_2_3_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_2_3_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_2_3_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_2_3_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_2_3_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_2_3_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_2_3_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_2_3_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_2_3_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_2_3_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_1_3_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_2_4_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_2_2_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_3_3_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_1_3_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_2_4_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_2_2_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_3_3_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_1_3_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_2_4_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_2_2_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_3_3_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_2_3_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_2_3_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_2_3_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_2_3_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_2_3_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_2_3_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_2_3_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_2_3_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_2_3_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_2_3_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_2_3_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_2_3_out_S_noc3_yummy )
);


tile
tile51 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[51] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd3),
    .default_coreid_y           (8'd3),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd51)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[51]   )
    ,.unavailable_o       ( unavailable_o[51] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[51]   )
    ,.ipi_i               ( ipi_i[51]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[51*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile51_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile51_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_2_3_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_3_4_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_3_2_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_4_3_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_2_3_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_3_4_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_3_2_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_4_3_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_2_3_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_3_4_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_3_2_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_4_3_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_3_3_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_3_3_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_3_3_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_3_3_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_3_3_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_3_3_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_3_3_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_3_3_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_3_3_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_3_3_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_3_3_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_3_3_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_2_3_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_3_4_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_3_2_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_4_3_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_2_3_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_3_4_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_3_2_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_4_3_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_2_3_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_3_4_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_3_2_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_4_3_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_3_3_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_3_3_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_3_3_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_3_3_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_3_3_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_3_3_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_3_3_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_3_3_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_3_3_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_3_3_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_3_3_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_3_3_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_2_3_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_3_4_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_3_2_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_4_3_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_2_3_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_3_4_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_3_2_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_4_3_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_2_3_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_3_4_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_3_2_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_4_3_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_3_3_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_3_3_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_3_3_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_3_3_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_3_3_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_3_3_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_3_3_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_3_3_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_3_3_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_3_3_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_3_3_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_3_3_out_S_noc3_yummy )
);


tile
tile67 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[67] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd3),
    .default_coreid_y           (8'd4),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd67)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[67]   )
    ,.unavailable_o       ( unavailable_o[67] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[67]   )
    ,.ipi_i               ( ipi_i[67]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[67*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile67_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile67_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_3_3_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_4_4_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_4_2_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_5_3_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_3_3_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_4_4_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_4_2_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_5_3_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_3_3_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_4_4_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_4_2_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_5_3_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_4_3_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_4_3_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_4_3_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_4_3_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_4_3_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_4_3_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_4_3_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_4_3_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_4_3_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_4_3_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_4_3_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_4_3_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_3_3_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_4_4_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_4_2_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_5_3_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_3_3_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_4_4_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_4_2_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_5_3_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_3_3_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_4_4_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_4_2_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_5_3_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_4_3_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_4_3_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_4_3_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_4_3_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_4_3_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_4_3_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_4_3_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_4_3_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_4_3_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_4_3_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_4_3_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_4_3_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_3_3_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_4_4_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_4_2_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_5_3_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_3_3_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_4_4_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_4_2_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_5_3_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_3_3_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_4_4_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_4_2_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_5_3_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_4_3_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_4_3_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_4_3_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_4_3_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_4_3_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_4_3_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_4_3_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_4_3_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_4_3_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_4_3_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_4_3_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_4_3_out_S_noc3_yummy )
);


tile
tile83 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[83] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd3),
    .default_coreid_y           (8'd5),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd83)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[83]   )
    ,.unavailable_o       ( unavailable_o[83] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[83]   )
    ,.ipi_i               ( ipi_i[83]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[83*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile83_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile83_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_4_3_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_5_4_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_5_2_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_6_3_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_4_3_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_5_4_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_5_2_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_6_3_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_4_3_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_5_4_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_5_2_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_6_3_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_5_3_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_5_3_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_5_3_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_5_3_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_5_3_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_5_3_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_5_3_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_5_3_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_5_3_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_5_3_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_5_3_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_5_3_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_4_3_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_5_4_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_5_2_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_6_3_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_4_3_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_5_4_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_5_2_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_6_3_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_4_3_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_5_4_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_5_2_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_6_3_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_5_3_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_5_3_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_5_3_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_5_3_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_5_3_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_5_3_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_5_3_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_5_3_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_5_3_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_5_3_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_5_3_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_5_3_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_4_3_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_5_4_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_5_2_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_6_3_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_4_3_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_5_4_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_5_2_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_6_3_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_4_3_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_5_4_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_5_2_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_6_3_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_5_3_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_5_3_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_5_3_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_5_3_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_5_3_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_5_3_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_5_3_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_5_3_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_5_3_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_5_3_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_5_3_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_5_3_out_S_noc3_yummy )
);


tile
tile99 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[99] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd3),
    .default_coreid_y           (8'd6),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd99)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[99]   )
    ,.unavailable_o       ( unavailable_o[99] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[99]   )
    ,.ipi_i               ( ipi_i[99]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[99*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile99_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile99_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_5_3_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_6_4_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_6_2_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_7_3_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_5_3_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_6_4_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_6_2_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_7_3_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_5_3_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_6_4_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_6_2_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_7_3_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_6_3_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_6_3_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_6_3_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_6_3_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_6_3_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_6_3_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_6_3_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_6_3_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_6_3_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_6_3_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_6_3_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_6_3_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_5_3_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_6_4_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_6_2_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_7_3_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_5_3_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_6_4_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_6_2_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_7_3_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_5_3_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_6_4_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_6_2_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_7_3_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_6_3_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_6_3_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_6_3_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_6_3_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_6_3_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_6_3_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_6_3_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_6_3_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_6_3_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_6_3_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_6_3_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_6_3_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_5_3_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_6_4_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_6_2_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_7_3_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_5_3_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_6_4_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_6_2_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_7_3_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_5_3_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_6_4_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_6_2_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_7_3_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_6_3_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_6_3_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_6_3_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_6_3_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_6_3_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_6_3_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_6_3_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_6_3_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_6_3_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_6_3_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_6_3_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_6_3_out_S_noc3_yummy )
);


tile
tile115 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[115] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd3),
    .default_coreid_y           (8'd7),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd115)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[115]   )
    ,.unavailable_o       ( unavailable_o[115] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[115]   )
    ,.ipi_i               ( ipi_i[115]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[115*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile115_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile115_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_6_3_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_7_4_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_7_2_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_8_3_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_6_3_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_7_4_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_7_2_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_8_3_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_6_3_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_7_4_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_7_2_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_8_3_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_7_3_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_7_3_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_7_3_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_7_3_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_7_3_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_7_3_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_7_3_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_7_3_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_7_3_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_7_3_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_7_3_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_7_3_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_6_3_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_7_4_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_7_2_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_8_3_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_6_3_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_7_4_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_7_2_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_8_3_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_6_3_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_7_4_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_7_2_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_8_3_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_7_3_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_7_3_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_7_3_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_7_3_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_7_3_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_7_3_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_7_3_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_7_3_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_7_3_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_7_3_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_7_3_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_7_3_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_6_3_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_7_4_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_7_2_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_8_3_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_6_3_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_7_4_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_7_2_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_8_3_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_6_3_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_7_4_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_7_2_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_8_3_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_7_3_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_7_3_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_7_3_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_7_3_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_7_3_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_7_3_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_7_3_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_7_3_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_7_3_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_7_3_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_7_3_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_7_3_out_S_noc3_yummy )
);


tile
tile131 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[131] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd3),
    .default_coreid_y           (8'd8),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd131)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[131]   )
    ,.unavailable_o       ( unavailable_o[131] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[131]   )
    ,.ipi_i               ( ipi_i[131]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[131*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile131_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile131_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_7_3_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_8_4_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_8_2_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_9_3_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_7_3_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_8_4_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_8_2_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_9_3_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_7_3_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_8_4_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_8_2_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_9_3_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_8_3_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_8_3_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_8_3_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_8_3_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_8_3_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_8_3_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_8_3_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_8_3_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_8_3_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_8_3_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_8_3_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_8_3_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_7_3_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_8_4_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_8_2_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_9_3_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_7_3_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_8_4_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_8_2_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_9_3_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_7_3_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_8_4_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_8_2_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_9_3_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_8_3_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_8_3_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_8_3_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_8_3_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_8_3_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_8_3_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_8_3_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_8_3_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_8_3_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_8_3_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_8_3_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_8_3_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_7_3_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_8_4_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_8_2_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_9_3_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_7_3_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_8_4_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_8_2_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_9_3_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_7_3_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_8_4_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_8_2_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_9_3_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_8_3_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_8_3_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_8_3_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_8_3_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_8_3_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_8_3_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_8_3_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_8_3_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_8_3_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_8_3_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_8_3_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_8_3_out_S_noc3_yummy )
);


tile
tile147 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[147] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd3),
    .default_coreid_y           (8'd9),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd147)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[147]   )
    ,.unavailable_o       ( unavailable_o[147] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[147]   )
    ,.ipi_i               ( ipi_i[147]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[147*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile147_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile147_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_8_3_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_9_4_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_9_2_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_10_3_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_8_3_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_9_4_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_9_2_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_10_3_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_8_3_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_9_4_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_9_2_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_10_3_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_9_3_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_9_3_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_9_3_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_9_3_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_9_3_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_9_3_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_9_3_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_9_3_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_9_3_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_9_3_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_9_3_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_9_3_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_8_3_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_9_4_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_9_2_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_10_3_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_8_3_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_9_4_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_9_2_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_10_3_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_8_3_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_9_4_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_9_2_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_10_3_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_9_3_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_9_3_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_9_3_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_9_3_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_9_3_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_9_3_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_9_3_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_9_3_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_9_3_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_9_3_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_9_3_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_9_3_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_8_3_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_9_4_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_9_2_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_10_3_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_8_3_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_9_4_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_9_2_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_10_3_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_8_3_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_9_4_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_9_2_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_10_3_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_9_3_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_9_3_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_9_3_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_9_3_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_9_3_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_9_3_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_9_3_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_9_3_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_9_3_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_9_3_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_9_3_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_9_3_out_S_noc3_yummy )
);


tile
tile163 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[163] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd3),
    .default_coreid_y           (8'd10),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd163)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[163]   )
    ,.unavailable_o       ( unavailable_o[163] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[163]   )
    ,.ipi_i               ( ipi_i[163]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[163*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile163_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile163_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_9_3_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_10_4_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_10_2_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_11_3_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_9_3_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_10_4_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_10_2_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_11_3_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_9_3_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_10_4_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_10_2_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_11_3_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_10_3_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_10_3_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_10_3_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_10_3_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_10_3_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_10_3_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_10_3_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_10_3_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_10_3_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_10_3_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_10_3_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_10_3_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_9_3_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_10_4_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_10_2_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_11_3_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_9_3_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_10_4_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_10_2_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_11_3_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_9_3_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_10_4_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_10_2_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_11_3_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_10_3_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_10_3_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_10_3_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_10_3_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_10_3_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_10_3_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_10_3_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_10_3_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_10_3_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_10_3_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_10_3_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_10_3_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_9_3_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_10_4_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_10_2_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_11_3_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_9_3_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_10_4_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_10_2_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_11_3_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_9_3_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_10_4_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_10_2_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_11_3_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_10_3_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_10_3_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_10_3_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_10_3_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_10_3_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_10_3_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_10_3_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_10_3_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_10_3_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_10_3_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_10_3_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_10_3_out_S_noc3_yummy )
);


tile
tile179 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[179] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd3),
    .default_coreid_y           (8'd11),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd179)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[179]   )
    ,.unavailable_o       ( unavailable_o[179] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[179]   )
    ,.ipi_i               ( ipi_i[179]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[179*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile179_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile179_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_10_3_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_11_4_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_11_2_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_12_3_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_10_3_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_11_4_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_11_2_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_12_3_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_10_3_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_11_4_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_11_2_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_12_3_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_11_3_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_11_3_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_11_3_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_11_3_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_11_3_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_11_3_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_11_3_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_11_3_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_11_3_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_11_3_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_11_3_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_11_3_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_10_3_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_11_4_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_11_2_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_12_3_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_10_3_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_11_4_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_11_2_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_12_3_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_10_3_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_11_4_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_11_2_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_12_3_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_11_3_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_11_3_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_11_3_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_11_3_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_11_3_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_11_3_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_11_3_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_11_3_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_11_3_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_11_3_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_11_3_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_11_3_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_10_3_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_11_4_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_11_2_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_12_3_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_10_3_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_11_4_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_11_2_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_12_3_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_10_3_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_11_4_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_11_2_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_12_3_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_11_3_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_11_3_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_11_3_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_11_3_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_11_3_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_11_3_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_11_3_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_11_3_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_11_3_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_11_3_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_11_3_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_11_3_out_S_noc3_yummy )
);


tile
tile195 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[195] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd3),
    .default_coreid_y           (8'd12),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd195)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[195]   )
    ,.unavailable_o       ( unavailable_o[195] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[195]   )
    ,.ipi_i               ( ipi_i[195]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[195*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile195_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile195_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_11_3_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_12_4_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_12_2_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_13_3_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_11_3_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_12_4_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_12_2_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_13_3_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_11_3_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_12_4_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_12_2_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_13_3_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_12_3_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_12_3_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_12_3_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_12_3_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_12_3_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_12_3_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_12_3_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_12_3_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_12_3_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_12_3_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_12_3_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_12_3_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_11_3_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_12_4_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_12_2_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_13_3_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_11_3_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_12_4_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_12_2_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_13_3_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_11_3_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_12_4_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_12_2_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_13_3_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_12_3_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_12_3_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_12_3_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_12_3_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_12_3_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_12_3_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_12_3_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_12_3_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_12_3_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_12_3_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_12_3_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_12_3_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_11_3_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_12_4_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_12_2_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_13_3_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_11_3_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_12_4_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_12_2_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_13_3_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_11_3_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_12_4_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_12_2_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_13_3_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_12_3_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_12_3_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_12_3_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_12_3_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_12_3_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_12_3_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_12_3_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_12_3_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_12_3_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_12_3_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_12_3_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_12_3_out_S_noc3_yummy )
);


tile
tile211 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[211] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd3),
    .default_coreid_y           (8'd13),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd211)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[211]   )
    ,.unavailable_o       ( unavailable_o[211] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[211]   )
    ,.ipi_i               ( ipi_i[211]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[211*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile211_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile211_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_12_3_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_13_4_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_13_2_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_14_3_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_12_3_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_13_4_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_13_2_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_14_3_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_12_3_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_13_4_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_13_2_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_14_3_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_13_3_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_13_3_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_13_3_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_13_3_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_13_3_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_13_3_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_13_3_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_13_3_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_13_3_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_13_3_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_13_3_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_13_3_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_12_3_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_13_4_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_13_2_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_14_3_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_12_3_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_13_4_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_13_2_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_14_3_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_12_3_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_13_4_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_13_2_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_14_3_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_13_3_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_13_3_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_13_3_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_13_3_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_13_3_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_13_3_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_13_3_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_13_3_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_13_3_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_13_3_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_13_3_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_13_3_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_12_3_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_13_4_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_13_2_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_14_3_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_12_3_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_13_4_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_13_2_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_14_3_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_12_3_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_13_4_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_13_2_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_14_3_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_13_3_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_13_3_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_13_3_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_13_3_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_13_3_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_13_3_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_13_3_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_13_3_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_13_3_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_13_3_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_13_3_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_13_3_out_S_noc3_yummy )
);


tile
tile227 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[227] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd3),
    .default_coreid_y           (8'd14),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd227)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[227]   )
    ,.unavailable_o       ( unavailable_o[227] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[227]   )
    ,.ipi_i               ( ipi_i[227]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[227*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile227_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile227_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_13_3_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_14_4_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_14_2_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_15_3_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_13_3_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_14_4_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_14_2_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_15_3_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_13_3_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_14_4_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_14_2_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_15_3_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_14_3_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_14_3_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_14_3_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_14_3_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_14_3_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_14_3_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_14_3_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_14_3_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_14_3_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_14_3_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_14_3_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_14_3_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_13_3_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_14_4_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_14_2_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_15_3_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_13_3_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_14_4_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_14_2_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_15_3_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_13_3_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_14_4_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_14_2_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_15_3_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_14_3_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_14_3_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_14_3_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_14_3_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_14_3_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_14_3_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_14_3_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_14_3_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_14_3_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_14_3_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_14_3_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_14_3_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_13_3_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_14_4_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_14_2_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_15_3_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_13_3_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_14_4_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_14_2_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_15_3_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_13_3_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_14_4_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_14_2_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_15_3_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_14_3_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_14_3_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_14_3_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_14_3_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_14_3_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_14_3_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_14_3_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_14_3_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_14_3_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_14_3_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_14_3_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_14_3_out_S_noc3_yummy )
);


tile
tile243 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[243] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd3),
    .default_coreid_y           (8'd15),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd243)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[243]   )
    ,.unavailable_o       ( unavailable_o[243] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[243]   )
    ,.ipi_i               ( ipi_i[243]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[243*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile243_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile243_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_14_3_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_15_4_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_15_2_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( dummy_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_14_3_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_15_4_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_15_2_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( dummy_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_14_3_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_15_4_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_15_2_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( dummy_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_15_3_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_15_3_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_15_3_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_15_3_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_15_3_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_15_3_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_15_3_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_15_3_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_15_3_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_15_3_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_15_3_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_15_3_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_14_3_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_15_4_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_15_2_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( dummy_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_14_3_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_15_4_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_15_2_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( dummy_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_14_3_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_15_4_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_15_2_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( dummy_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_15_3_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_15_3_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_15_3_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_15_3_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_15_3_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_15_3_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_15_3_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_15_3_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_15_3_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_15_3_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_15_3_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_15_3_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_14_3_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_15_4_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_15_2_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( dummy_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_14_3_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_15_4_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_15_2_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( dummy_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_14_3_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_15_4_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_15_2_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( dummy_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_15_3_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_15_3_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_15_3_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_15_3_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_15_3_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_15_3_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_15_3_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_15_3_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_15_3_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_15_3_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_15_3_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_15_3_out_S_noc3_yummy )
);


tile
tile4 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[4] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd4),
    .default_coreid_y           (8'd0),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd4)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[4]   )
    ,.unavailable_o       ( unavailable_o[4] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[4]   )
    ,.ipi_i               ( ipi_i[4]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[4*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile4_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile4_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( dummy_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_0_5_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_0_3_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_1_4_out_N_noc1_data   ),
    .dyn0_validIn_N      ( dummy_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_0_5_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_0_3_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_1_4_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( dummy_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_0_5_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_0_3_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_1_4_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_0_4_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_0_4_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_0_4_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_0_4_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_0_4_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_0_4_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_0_4_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_0_4_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_0_4_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_0_4_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_0_4_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_0_4_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( dummy_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_0_5_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_0_3_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_1_4_out_N_noc2_data   ),
    .dyn1_validIn_N      ( dummy_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_0_5_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_0_3_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_1_4_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( dummy_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_0_5_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_0_3_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_1_4_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_0_4_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_0_4_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_0_4_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_0_4_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_0_4_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_0_4_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_0_4_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_0_4_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_0_4_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_0_4_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_0_4_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_0_4_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( dummy_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_0_5_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_0_3_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_1_4_out_N_noc3_data   ),
    .dyn2_validIn_N      ( dummy_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_0_5_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_0_3_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_1_4_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( dummy_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_0_5_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_0_3_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_1_4_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_0_4_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_0_4_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_0_4_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_0_4_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_0_4_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_0_4_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_0_4_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_0_4_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_0_4_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_0_4_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_0_4_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_0_4_out_S_noc3_yummy )
);


tile
tile20 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[20] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd4),
    .default_coreid_y           (8'd1),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd20)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[20]   )
    ,.unavailable_o       ( unavailable_o[20] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[20]   )
    ,.ipi_i               ( ipi_i[20]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[20*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile20_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile20_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_0_4_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_1_5_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_1_3_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_2_4_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_0_4_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_1_5_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_1_3_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_2_4_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_0_4_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_1_5_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_1_3_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_2_4_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_1_4_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_1_4_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_1_4_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_1_4_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_1_4_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_1_4_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_1_4_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_1_4_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_1_4_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_1_4_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_1_4_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_1_4_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_0_4_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_1_5_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_1_3_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_2_4_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_0_4_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_1_5_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_1_3_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_2_4_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_0_4_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_1_5_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_1_3_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_2_4_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_1_4_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_1_4_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_1_4_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_1_4_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_1_4_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_1_4_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_1_4_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_1_4_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_1_4_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_1_4_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_1_4_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_1_4_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_0_4_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_1_5_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_1_3_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_2_4_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_0_4_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_1_5_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_1_3_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_2_4_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_0_4_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_1_5_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_1_3_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_2_4_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_1_4_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_1_4_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_1_4_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_1_4_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_1_4_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_1_4_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_1_4_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_1_4_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_1_4_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_1_4_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_1_4_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_1_4_out_S_noc3_yummy )
);


tile
tile36 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[36] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd4),
    .default_coreid_y           (8'd2),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd36)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[36]   )
    ,.unavailable_o       ( unavailable_o[36] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[36]   )
    ,.ipi_i               ( ipi_i[36]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[36*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile36_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile36_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_1_4_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_2_5_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_2_3_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_3_4_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_1_4_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_2_5_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_2_3_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_3_4_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_1_4_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_2_5_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_2_3_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_3_4_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_2_4_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_2_4_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_2_4_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_2_4_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_2_4_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_2_4_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_2_4_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_2_4_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_2_4_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_2_4_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_2_4_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_2_4_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_1_4_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_2_5_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_2_3_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_3_4_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_1_4_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_2_5_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_2_3_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_3_4_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_1_4_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_2_5_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_2_3_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_3_4_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_2_4_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_2_4_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_2_4_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_2_4_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_2_4_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_2_4_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_2_4_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_2_4_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_2_4_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_2_4_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_2_4_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_2_4_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_1_4_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_2_5_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_2_3_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_3_4_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_1_4_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_2_5_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_2_3_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_3_4_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_1_4_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_2_5_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_2_3_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_3_4_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_2_4_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_2_4_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_2_4_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_2_4_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_2_4_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_2_4_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_2_4_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_2_4_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_2_4_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_2_4_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_2_4_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_2_4_out_S_noc3_yummy )
);


tile
tile52 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[52] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd4),
    .default_coreid_y           (8'd3),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd52)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[52]   )
    ,.unavailable_o       ( unavailable_o[52] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[52]   )
    ,.ipi_i               ( ipi_i[52]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[52*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile52_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile52_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_2_4_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_3_5_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_3_3_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_4_4_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_2_4_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_3_5_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_3_3_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_4_4_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_2_4_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_3_5_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_3_3_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_4_4_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_3_4_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_3_4_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_3_4_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_3_4_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_3_4_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_3_4_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_3_4_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_3_4_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_3_4_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_3_4_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_3_4_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_3_4_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_2_4_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_3_5_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_3_3_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_4_4_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_2_4_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_3_5_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_3_3_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_4_4_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_2_4_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_3_5_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_3_3_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_4_4_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_3_4_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_3_4_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_3_4_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_3_4_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_3_4_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_3_4_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_3_4_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_3_4_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_3_4_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_3_4_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_3_4_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_3_4_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_2_4_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_3_5_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_3_3_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_4_4_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_2_4_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_3_5_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_3_3_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_4_4_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_2_4_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_3_5_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_3_3_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_4_4_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_3_4_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_3_4_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_3_4_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_3_4_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_3_4_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_3_4_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_3_4_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_3_4_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_3_4_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_3_4_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_3_4_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_3_4_out_S_noc3_yummy )
);


tile
tile68 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[68] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd4),
    .default_coreid_y           (8'd4),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd68)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[68]   )
    ,.unavailable_o       ( unavailable_o[68] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[68]   )
    ,.ipi_i               ( ipi_i[68]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[68*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile68_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile68_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_3_4_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_4_5_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_4_3_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_5_4_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_3_4_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_4_5_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_4_3_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_5_4_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_3_4_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_4_5_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_4_3_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_5_4_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_4_4_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_4_4_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_4_4_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_4_4_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_4_4_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_4_4_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_4_4_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_4_4_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_4_4_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_4_4_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_4_4_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_4_4_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_3_4_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_4_5_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_4_3_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_5_4_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_3_4_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_4_5_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_4_3_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_5_4_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_3_4_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_4_5_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_4_3_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_5_4_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_4_4_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_4_4_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_4_4_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_4_4_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_4_4_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_4_4_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_4_4_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_4_4_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_4_4_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_4_4_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_4_4_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_4_4_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_3_4_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_4_5_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_4_3_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_5_4_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_3_4_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_4_5_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_4_3_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_5_4_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_3_4_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_4_5_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_4_3_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_5_4_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_4_4_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_4_4_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_4_4_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_4_4_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_4_4_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_4_4_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_4_4_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_4_4_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_4_4_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_4_4_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_4_4_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_4_4_out_S_noc3_yummy )
);


tile
tile84 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[84] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd4),
    .default_coreid_y           (8'd5),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd84)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[84]   )
    ,.unavailable_o       ( unavailable_o[84] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[84]   )
    ,.ipi_i               ( ipi_i[84]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[84*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile84_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile84_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_4_4_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_5_5_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_5_3_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_6_4_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_4_4_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_5_5_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_5_3_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_6_4_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_4_4_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_5_5_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_5_3_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_6_4_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_5_4_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_5_4_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_5_4_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_5_4_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_5_4_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_5_4_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_5_4_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_5_4_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_5_4_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_5_4_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_5_4_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_5_4_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_4_4_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_5_5_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_5_3_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_6_4_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_4_4_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_5_5_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_5_3_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_6_4_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_4_4_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_5_5_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_5_3_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_6_4_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_5_4_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_5_4_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_5_4_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_5_4_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_5_4_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_5_4_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_5_4_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_5_4_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_5_4_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_5_4_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_5_4_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_5_4_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_4_4_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_5_5_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_5_3_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_6_4_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_4_4_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_5_5_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_5_3_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_6_4_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_4_4_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_5_5_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_5_3_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_6_4_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_5_4_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_5_4_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_5_4_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_5_4_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_5_4_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_5_4_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_5_4_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_5_4_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_5_4_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_5_4_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_5_4_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_5_4_out_S_noc3_yummy )
);


tile
tile100 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[100] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd4),
    .default_coreid_y           (8'd6),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd100)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[100]   )
    ,.unavailable_o       ( unavailable_o[100] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[100]   )
    ,.ipi_i               ( ipi_i[100]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[100*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile100_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile100_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_5_4_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_6_5_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_6_3_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_7_4_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_5_4_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_6_5_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_6_3_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_7_4_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_5_4_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_6_5_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_6_3_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_7_4_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_6_4_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_6_4_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_6_4_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_6_4_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_6_4_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_6_4_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_6_4_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_6_4_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_6_4_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_6_4_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_6_4_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_6_4_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_5_4_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_6_5_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_6_3_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_7_4_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_5_4_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_6_5_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_6_3_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_7_4_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_5_4_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_6_5_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_6_3_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_7_4_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_6_4_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_6_4_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_6_4_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_6_4_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_6_4_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_6_4_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_6_4_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_6_4_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_6_4_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_6_4_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_6_4_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_6_4_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_5_4_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_6_5_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_6_3_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_7_4_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_5_4_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_6_5_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_6_3_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_7_4_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_5_4_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_6_5_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_6_3_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_7_4_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_6_4_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_6_4_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_6_4_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_6_4_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_6_4_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_6_4_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_6_4_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_6_4_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_6_4_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_6_4_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_6_4_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_6_4_out_S_noc3_yummy )
);


tile
tile116 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[116] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd4),
    .default_coreid_y           (8'd7),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd116)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[116]   )
    ,.unavailable_o       ( unavailable_o[116] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[116]   )
    ,.ipi_i               ( ipi_i[116]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[116*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile116_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile116_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_6_4_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_7_5_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_7_3_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_8_4_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_6_4_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_7_5_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_7_3_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_8_4_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_6_4_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_7_5_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_7_3_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_8_4_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_7_4_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_7_4_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_7_4_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_7_4_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_7_4_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_7_4_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_7_4_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_7_4_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_7_4_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_7_4_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_7_4_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_7_4_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_6_4_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_7_5_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_7_3_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_8_4_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_6_4_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_7_5_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_7_3_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_8_4_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_6_4_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_7_5_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_7_3_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_8_4_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_7_4_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_7_4_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_7_4_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_7_4_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_7_4_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_7_4_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_7_4_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_7_4_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_7_4_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_7_4_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_7_4_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_7_4_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_6_4_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_7_5_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_7_3_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_8_4_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_6_4_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_7_5_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_7_3_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_8_4_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_6_4_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_7_5_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_7_3_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_8_4_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_7_4_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_7_4_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_7_4_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_7_4_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_7_4_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_7_4_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_7_4_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_7_4_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_7_4_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_7_4_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_7_4_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_7_4_out_S_noc3_yummy )
);


tile
tile132 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[132] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd4),
    .default_coreid_y           (8'd8),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd132)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[132]   )
    ,.unavailable_o       ( unavailable_o[132] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[132]   )
    ,.ipi_i               ( ipi_i[132]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[132*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile132_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile132_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_7_4_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_8_5_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_8_3_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_9_4_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_7_4_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_8_5_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_8_3_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_9_4_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_7_4_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_8_5_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_8_3_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_9_4_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_8_4_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_8_4_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_8_4_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_8_4_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_8_4_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_8_4_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_8_4_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_8_4_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_8_4_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_8_4_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_8_4_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_8_4_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_7_4_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_8_5_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_8_3_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_9_4_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_7_4_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_8_5_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_8_3_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_9_4_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_7_4_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_8_5_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_8_3_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_9_4_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_8_4_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_8_4_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_8_4_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_8_4_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_8_4_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_8_4_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_8_4_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_8_4_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_8_4_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_8_4_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_8_4_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_8_4_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_7_4_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_8_5_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_8_3_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_9_4_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_7_4_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_8_5_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_8_3_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_9_4_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_7_4_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_8_5_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_8_3_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_9_4_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_8_4_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_8_4_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_8_4_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_8_4_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_8_4_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_8_4_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_8_4_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_8_4_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_8_4_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_8_4_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_8_4_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_8_4_out_S_noc3_yummy )
);


tile
tile148 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[148] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd4),
    .default_coreid_y           (8'd9),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd148)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[148]   )
    ,.unavailable_o       ( unavailable_o[148] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[148]   )
    ,.ipi_i               ( ipi_i[148]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[148*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile148_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile148_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_8_4_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_9_5_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_9_3_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_10_4_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_8_4_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_9_5_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_9_3_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_10_4_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_8_4_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_9_5_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_9_3_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_10_4_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_9_4_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_9_4_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_9_4_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_9_4_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_9_4_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_9_4_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_9_4_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_9_4_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_9_4_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_9_4_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_9_4_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_9_4_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_8_4_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_9_5_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_9_3_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_10_4_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_8_4_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_9_5_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_9_3_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_10_4_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_8_4_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_9_5_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_9_3_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_10_4_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_9_4_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_9_4_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_9_4_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_9_4_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_9_4_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_9_4_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_9_4_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_9_4_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_9_4_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_9_4_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_9_4_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_9_4_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_8_4_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_9_5_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_9_3_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_10_4_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_8_4_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_9_5_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_9_3_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_10_4_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_8_4_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_9_5_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_9_3_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_10_4_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_9_4_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_9_4_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_9_4_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_9_4_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_9_4_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_9_4_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_9_4_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_9_4_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_9_4_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_9_4_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_9_4_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_9_4_out_S_noc3_yummy )
);


tile
tile164 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[164] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd4),
    .default_coreid_y           (8'd10),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd164)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[164]   )
    ,.unavailable_o       ( unavailable_o[164] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[164]   )
    ,.ipi_i               ( ipi_i[164]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[164*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile164_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile164_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_9_4_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_10_5_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_10_3_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_11_4_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_9_4_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_10_5_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_10_3_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_11_4_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_9_4_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_10_5_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_10_3_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_11_4_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_10_4_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_10_4_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_10_4_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_10_4_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_10_4_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_10_4_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_10_4_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_10_4_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_10_4_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_10_4_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_10_4_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_10_4_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_9_4_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_10_5_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_10_3_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_11_4_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_9_4_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_10_5_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_10_3_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_11_4_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_9_4_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_10_5_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_10_3_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_11_4_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_10_4_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_10_4_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_10_4_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_10_4_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_10_4_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_10_4_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_10_4_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_10_4_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_10_4_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_10_4_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_10_4_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_10_4_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_9_4_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_10_5_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_10_3_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_11_4_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_9_4_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_10_5_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_10_3_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_11_4_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_9_4_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_10_5_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_10_3_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_11_4_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_10_4_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_10_4_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_10_4_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_10_4_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_10_4_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_10_4_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_10_4_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_10_4_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_10_4_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_10_4_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_10_4_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_10_4_out_S_noc3_yummy )
);


tile
tile180 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[180] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd4),
    .default_coreid_y           (8'd11),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd180)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[180]   )
    ,.unavailable_o       ( unavailable_o[180] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[180]   )
    ,.ipi_i               ( ipi_i[180]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[180*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile180_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile180_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_10_4_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_11_5_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_11_3_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_12_4_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_10_4_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_11_5_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_11_3_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_12_4_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_10_4_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_11_5_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_11_3_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_12_4_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_11_4_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_11_4_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_11_4_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_11_4_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_11_4_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_11_4_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_11_4_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_11_4_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_11_4_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_11_4_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_11_4_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_11_4_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_10_4_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_11_5_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_11_3_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_12_4_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_10_4_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_11_5_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_11_3_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_12_4_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_10_4_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_11_5_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_11_3_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_12_4_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_11_4_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_11_4_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_11_4_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_11_4_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_11_4_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_11_4_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_11_4_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_11_4_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_11_4_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_11_4_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_11_4_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_11_4_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_10_4_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_11_5_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_11_3_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_12_4_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_10_4_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_11_5_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_11_3_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_12_4_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_10_4_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_11_5_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_11_3_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_12_4_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_11_4_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_11_4_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_11_4_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_11_4_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_11_4_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_11_4_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_11_4_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_11_4_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_11_4_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_11_4_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_11_4_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_11_4_out_S_noc3_yummy )
);


tile
tile196 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[196] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd4),
    .default_coreid_y           (8'd12),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd196)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[196]   )
    ,.unavailable_o       ( unavailable_o[196] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[196]   )
    ,.ipi_i               ( ipi_i[196]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[196*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile196_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile196_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_11_4_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_12_5_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_12_3_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_13_4_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_11_4_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_12_5_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_12_3_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_13_4_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_11_4_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_12_5_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_12_3_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_13_4_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_12_4_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_12_4_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_12_4_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_12_4_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_12_4_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_12_4_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_12_4_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_12_4_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_12_4_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_12_4_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_12_4_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_12_4_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_11_4_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_12_5_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_12_3_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_13_4_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_11_4_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_12_5_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_12_3_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_13_4_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_11_4_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_12_5_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_12_3_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_13_4_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_12_4_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_12_4_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_12_4_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_12_4_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_12_4_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_12_4_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_12_4_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_12_4_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_12_4_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_12_4_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_12_4_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_12_4_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_11_4_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_12_5_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_12_3_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_13_4_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_11_4_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_12_5_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_12_3_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_13_4_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_11_4_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_12_5_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_12_3_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_13_4_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_12_4_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_12_4_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_12_4_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_12_4_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_12_4_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_12_4_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_12_4_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_12_4_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_12_4_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_12_4_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_12_4_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_12_4_out_S_noc3_yummy )
);


tile
tile212 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[212] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd4),
    .default_coreid_y           (8'd13),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd212)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[212]   )
    ,.unavailable_o       ( unavailable_o[212] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[212]   )
    ,.ipi_i               ( ipi_i[212]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[212*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile212_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile212_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_12_4_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_13_5_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_13_3_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_14_4_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_12_4_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_13_5_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_13_3_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_14_4_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_12_4_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_13_5_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_13_3_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_14_4_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_13_4_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_13_4_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_13_4_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_13_4_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_13_4_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_13_4_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_13_4_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_13_4_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_13_4_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_13_4_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_13_4_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_13_4_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_12_4_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_13_5_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_13_3_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_14_4_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_12_4_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_13_5_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_13_3_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_14_4_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_12_4_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_13_5_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_13_3_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_14_4_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_13_4_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_13_4_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_13_4_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_13_4_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_13_4_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_13_4_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_13_4_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_13_4_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_13_4_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_13_4_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_13_4_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_13_4_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_12_4_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_13_5_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_13_3_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_14_4_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_12_4_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_13_5_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_13_3_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_14_4_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_12_4_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_13_5_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_13_3_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_14_4_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_13_4_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_13_4_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_13_4_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_13_4_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_13_4_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_13_4_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_13_4_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_13_4_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_13_4_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_13_4_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_13_4_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_13_4_out_S_noc3_yummy )
);


tile
tile228 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[228] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd4),
    .default_coreid_y           (8'd14),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd228)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[228]   )
    ,.unavailable_o       ( unavailable_o[228] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[228]   )
    ,.ipi_i               ( ipi_i[228]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[228*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile228_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile228_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_13_4_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_14_5_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_14_3_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_15_4_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_13_4_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_14_5_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_14_3_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_15_4_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_13_4_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_14_5_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_14_3_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_15_4_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_14_4_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_14_4_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_14_4_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_14_4_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_14_4_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_14_4_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_14_4_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_14_4_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_14_4_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_14_4_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_14_4_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_14_4_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_13_4_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_14_5_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_14_3_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_15_4_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_13_4_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_14_5_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_14_3_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_15_4_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_13_4_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_14_5_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_14_3_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_15_4_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_14_4_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_14_4_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_14_4_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_14_4_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_14_4_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_14_4_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_14_4_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_14_4_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_14_4_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_14_4_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_14_4_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_14_4_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_13_4_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_14_5_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_14_3_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_15_4_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_13_4_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_14_5_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_14_3_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_15_4_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_13_4_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_14_5_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_14_3_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_15_4_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_14_4_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_14_4_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_14_4_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_14_4_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_14_4_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_14_4_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_14_4_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_14_4_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_14_4_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_14_4_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_14_4_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_14_4_out_S_noc3_yummy )
);


tile
tile244 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[244] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd4),
    .default_coreid_y           (8'd15),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd244)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[244]   )
    ,.unavailable_o       ( unavailable_o[244] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[244]   )
    ,.ipi_i               ( ipi_i[244]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[244*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile244_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile244_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_14_4_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_15_5_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_15_3_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( dummy_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_14_4_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_15_5_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_15_3_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( dummy_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_14_4_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_15_5_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_15_3_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( dummy_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_15_4_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_15_4_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_15_4_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_15_4_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_15_4_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_15_4_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_15_4_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_15_4_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_15_4_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_15_4_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_15_4_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_15_4_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_14_4_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_15_5_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_15_3_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( dummy_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_14_4_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_15_5_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_15_3_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( dummy_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_14_4_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_15_5_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_15_3_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( dummy_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_15_4_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_15_4_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_15_4_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_15_4_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_15_4_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_15_4_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_15_4_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_15_4_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_15_4_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_15_4_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_15_4_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_15_4_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_14_4_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_15_5_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_15_3_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( dummy_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_14_4_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_15_5_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_15_3_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( dummy_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_14_4_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_15_5_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_15_3_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( dummy_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_15_4_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_15_4_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_15_4_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_15_4_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_15_4_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_15_4_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_15_4_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_15_4_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_15_4_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_15_4_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_15_4_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_15_4_out_S_noc3_yummy )
);


tile
tile5 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[5] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd5),
    .default_coreid_y           (8'd0),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd5)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[5]   )
    ,.unavailable_o       ( unavailable_o[5] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[5]   )
    ,.ipi_i               ( ipi_i[5]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[5*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile5_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile5_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( dummy_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_0_6_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_0_4_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_1_5_out_N_noc1_data   ),
    .dyn0_validIn_N      ( dummy_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_0_6_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_0_4_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_1_5_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( dummy_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_0_6_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_0_4_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_1_5_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_0_5_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_0_5_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_0_5_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_0_5_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_0_5_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_0_5_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_0_5_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_0_5_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_0_5_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_0_5_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_0_5_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_0_5_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( dummy_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_0_6_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_0_4_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_1_5_out_N_noc2_data   ),
    .dyn1_validIn_N      ( dummy_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_0_6_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_0_4_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_1_5_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( dummy_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_0_6_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_0_4_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_1_5_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_0_5_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_0_5_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_0_5_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_0_5_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_0_5_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_0_5_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_0_5_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_0_5_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_0_5_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_0_5_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_0_5_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_0_5_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( dummy_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_0_6_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_0_4_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_1_5_out_N_noc3_data   ),
    .dyn2_validIn_N      ( dummy_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_0_6_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_0_4_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_1_5_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( dummy_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_0_6_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_0_4_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_1_5_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_0_5_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_0_5_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_0_5_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_0_5_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_0_5_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_0_5_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_0_5_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_0_5_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_0_5_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_0_5_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_0_5_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_0_5_out_S_noc3_yummy )
);


tile
tile21 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[21] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd5),
    .default_coreid_y           (8'd1),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd21)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[21]   )
    ,.unavailable_o       ( unavailable_o[21] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[21]   )
    ,.ipi_i               ( ipi_i[21]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[21*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile21_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile21_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_0_5_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_1_6_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_1_4_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_2_5_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_0_5_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_1_6_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_1_4_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_2_5_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_0_5_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_1_6_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_1_4_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_2_5_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_1_5_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_1_5_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_1_5_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_1_5_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_1_5_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_1_5_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_1_5_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_1_5_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_1_5_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_1_5_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_1_5_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_1_5_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_0_5_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_1_6_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_1_4_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_2_5_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_0_5_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_1_6_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_1_4_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_2_5_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_0_5_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_1_6_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_1_4_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_2_5_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_1_5_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_1_5_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_1_5_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_1_5_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_1_5_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_1_5_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_1_5_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_1_5_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_1_5_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_1_5_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_1_5_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_1_5_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_0_5_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_1_6_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_1_4_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_2_5_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_0_5_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_1_6_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_1_4_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_2_5_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_0_5_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_1_6_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_1_4_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_2_5_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_1_5_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_1_5_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_1_5_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_1_5_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_1_5_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_1_5_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_1_5_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_1_5_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_1_5_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_1_5_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_1_5_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_1_5_out_S_noc3_yummy )
);


tile
tile37 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[37] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd5),
    .default_coreid_y           (8'd2),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd37)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[37]   )
    ,.unavailable_o       ( unavailable_o[37] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[37]   )
    ,.ipi_i               ( ipi_i[37]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[37*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile37_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile37_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_1_5_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_2_6_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_2_4_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_3_5_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_1_5_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_2_6_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_2_4_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_3_5_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_1_5_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_2_6_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_2_4_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_3_5_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_2_5_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_2_5_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_2_5_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_2_5_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_2_5_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_2_5_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_2_5_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_2_5_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_2_5_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_2_5_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_2_5_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_2_5_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_1_5_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_2_6_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_2_4_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_3_5_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_1_5_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_2_6_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_2_4_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_3_5_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_1_5_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_2_6_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_2_4_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_3_5_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_2_5_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_2_5_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_2_5_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_2_5_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_2_5_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_2_5_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_2_5_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_2_5_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_2_5_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_2_5_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_2_5_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_2_5_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_1_5_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_2_6_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_2_4_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_3_5_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_1_5_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_2_6_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_2_4_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_3_5_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_1_5_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_2_6_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_2_4_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_3_5_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_2_5_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_2_5_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_2_5_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_2_5_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_2_5_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_2_5_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_2_5_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_2_5_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_2_5_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_2_5_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_2_5_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_2_5_out_S_noc3_yummy )
);


tile
tile53 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[53] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd5),
    .default_coreid_y           (8'd3),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd53)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[53]   )
    ,.unavailable_o       ( unavailable_o[53] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[53]   )
    ,.ipi_i               ( ipi_i[53]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[53*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile53_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile53_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_2_5_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_3_6_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_3_4_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_4_5_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_2_5_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_3_6_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_3_4_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_4_5_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_2_5_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_3_6_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_3_4_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_4_5_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_3_5_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_3_5_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_3_5_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_3_5_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_3_5_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_3_5_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_3_5_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_3_5_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_3_5_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_3_5_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_3_5_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_3_5_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_2_5_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_3_6_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_3_4_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_4_5_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_2_5_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_3_6_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_3_4_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_4_5_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_2_5_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_3_6_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_3_4_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_4_5_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_3_5_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_3_5_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_3_5_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_3_5_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_3_5_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_3_5_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_3_5_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_3_5_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_3_5_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_3_5_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_3_5_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_3_5_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_2_5_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_3_6_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_3_4_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_4_5_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_2_5_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_3_6_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_3_4_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_4_5_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_2_5_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_3_6_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_3_4_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_4_5_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_3_5_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_3_5_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_3_5_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_3_5_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_3_5_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_3_5_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_3_5_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_3_5_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_3_5_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_3_5_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_3_5_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_3_5_out_S_noc3_yummy )
);


tile
tile69 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[69] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd5),
    .default_coreid_y           (8'd4),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd69)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[69]   )
    ,.unavailable_o       ( unavailable_o[69] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[69]   )
    ,.ipi_i               ( ipi_i[69]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[69*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile69_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile69_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_3_5_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_4_6_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_4_4_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_5_5_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_3_5_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_4_6_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_4_4_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_5_5_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_3_5_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_4_6_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_4_4_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_5_5_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_4_5_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_4_5_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_4_5_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_4_5_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_4_5_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_4_5_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_4_5_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_4_5_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_4_5_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_4_5_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_4_5_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_4_5_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_3_5_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_4_6_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_4_4_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_5_5_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_3_5_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_4_6_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_4_4_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_5_5_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_3_5_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_4_6_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_4_4_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_5_5_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_4_5_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_4_5_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_4_5_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_4_5_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_4_5_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_4_5_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_4_5_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_4_5_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_4_5_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_4_5_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_4_5_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_4_5_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_3_5_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_4_6_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_4_4_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_5_5_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_3_5_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_4_6_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_4_4_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_5_5_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_3_5_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_4_6_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_4_4_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_5_5_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_4_5_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_4_5_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_4_5_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_4_5_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_4_5_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_4_5_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_4_5_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_4_5_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_4_5_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_4_5_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_4_5_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_4_5_out_S_noc3_yummy )
);


tile
tile85 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[85] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd5),
    .default_coreid_y           (8'd5),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd85)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[85]   )
    ,.unavailable_o       ( unavailable_o[85] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[85]   )
    ,.ipi_i               ( ipi_i[85]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[85*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile85_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile85_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_4_5_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_5_6_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_5_4_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_6_5_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_4_5_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_5_6_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_5_4_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_6_5_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_4_5_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_5_6_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_5_4_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_6_5_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_5_5_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_5_5_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_5_5_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_5_5_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_5_5_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_5_5_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_5_5_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_5_5_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_5_5_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_5_5_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_5_5_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_5_5_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_4_5_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_5_6_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_5_4_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_6_5_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_4_5_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_5_6_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_5_4_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_6_5_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_4_5_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_5_6_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_5_4_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_6_5_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_5_5_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_5_5_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_5_5_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_5_5_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_5_5_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_5_5_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_5_5_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_5_5_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_5_5_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_5_5_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_5_5_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_5_5_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_4_5_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_5_6_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_5_4_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_6_5_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_4_5_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_5_6_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_5_4_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_6_5_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_4_5_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_5_6_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_5_4_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_6_5_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_5_5_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_5_5_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_5_5_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_5_5_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_5_5_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_5_5_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_5_5_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_5_5_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_5_5_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_5_5_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_5_5_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_5_5_out_S_noc3_yummy )
);


tile
tile101 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[101] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd5),
    .default_coreid_y           (8'd6),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd101)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[101]   )
    ,.unavailable_o       ( unavailable_o[101] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[101]   )
    ,.ipi_i               ( ipi_i[101]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[101*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile101_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile101_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_5_5_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_6_6_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_6_4_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_7_5_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_5_5_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_6_6_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_6_4_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_7_5_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_5_5_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_6_6_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_6_4_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_7_5_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_6_5_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_6_5_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_6_5_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_6_5_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_6_5_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_6_5_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_6_5_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_6_5_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_6_5_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_6_5_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_6_5_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_6_5_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_5_5_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_6_6_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_6_4_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_7_5_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_5_5_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_6_6_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_6_4_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_7_5_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_5_5_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_6_6_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_6_4_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_7_5_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_6_5_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_6_5_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_6_5_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_6_5_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_6_5_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_6_5_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_6_5_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_6_5_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_6_5_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_6_5_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_6_5_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_6_5_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_5_5_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_6_6_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_6_4_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_7_5_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_5_5_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_6_6_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_6_4_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_7_5_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_5_5_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_6_6_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_6_4_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_7_5_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_6_5_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_6_5_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_6_5_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_6_5_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_6_5_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_6_5_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_6_5_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_6_5_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_6_5_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_6_5_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_6_5_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_6_5_out_S_noc3_yummy )
);


tile
tile117 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[117] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd5),
    .default_coreid_y           (8'd7),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd117)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[117]   )
    ,.unavailable_o       ( unavailable_o[117] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[117]   )
    ,.ipi_i               ( ipi_i[117]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[117*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile117_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile117_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_6_5_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_7_6_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_7_4_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_8_5_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_6_5_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_7_6_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_7_4_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_8_5_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_6_5_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_7_6_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_7_4_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_8_5_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_7_5_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_7_5_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_7_5_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_7_5_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_7_5_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_7_5_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_7_5_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_7_5_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_7_5_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_7_5_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_7_5_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_7_5_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_6_5_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_7_6_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_7_4_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_8_5_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_6_5_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_7_6_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_7_4_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_8_5_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_6_5_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_7_6_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_7_4_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_8_5_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_7_5_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_7_5_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_7_5_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_7_5_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_7_5_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_7_5_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_7_5_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_7_5_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_7_5_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_7_5_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_7_5_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_7_5_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_6_5_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_7_6_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_7_4_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_8_5_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_6_5_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_7_6_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_7_4_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_8_5_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_6_5_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_7_6_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_7_4_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_8_5_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_7_5_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_7_5_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_7_5_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_7_5_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_7_5_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_7_5_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_7_5_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_7_5_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_7_5_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_7_5_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_7_5_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_7_5_out_S_noc3_yummy )
);


tile
tile133 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[133] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd5),
    .default_coreid_y           (8'd8),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd133)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[133]   )
    ,.unavailable_o       ( unavailable_o[133] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[133]   )
    ,.ipi_i               ( ipi_i[133]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[133*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile133_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile133_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_7_5_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_8_6_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_8_4_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_9_5_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_7_5_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_8_6_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_8_4_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_9_5_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_7_5_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_8_6_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_8_4_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_9_5_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_8_5_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_8_5_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_8_5_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_8_5_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_8_5_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_8_5_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_8_5_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_8_5_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_8_5_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_8_5_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_8_5_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_8_5_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_7_5_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_8_6_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_8_4_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_9_5_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_7_5_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_8_6_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_8_4_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_9_5_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_7_5_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_8_6_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_8_4_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_9_5_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_8_5_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_8_5_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_8_5_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_8_5_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_8_5_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_8_5_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_8_5_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_8_5_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_8_5_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_8_5_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_8_5_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_8_5_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_7_5_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_8_6_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_8_4_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_9_5_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_7_5_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_8_6_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_8_4_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_9_5_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_7_5_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_8_6_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_8_4_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_9_5_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_8_5_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_8_5_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_8_5_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_8_5_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_8_5_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_8_5_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_8_5_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_8_5_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_8_5_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_8_5_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_8_5_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_8_5_out_S_noc3_yummy )
);


tile
tile149 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[149] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd5),
    .default_coreid_y           (8'd9),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd149)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[149]   )
    ,.unavailable_o       ( unavailable_o[149] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[149]   )
    ,.ipi_i               ( ipi_i[149]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[149*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile149_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile149_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_8_5_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_9_6_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_9_4_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_10_5_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_8_5_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_9_6_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_9_4_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_10_5_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_8_5_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_9_6_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_9_4_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_10_5_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_9_5_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_9_5_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_9_5_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_9_5_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_9_5_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_9_5_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_9_5_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_9_5_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_9_5_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_9_5_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_9_5_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_9_5_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_8_5_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_9_6_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_9_4_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_10_5_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_8_5_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_9_6_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_9_4_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_10_5_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_8_5_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_9_6_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_9_4_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_10_5_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_9_5_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_9_5_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_9_5_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_9_5_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_9_5_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_9_5_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_9_5_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_9_5_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_9_5_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_9_5_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_9_5_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_9_5_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_8_5_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_9_6_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_9_4_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_10_5_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_8_5_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_9_6_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_9_4_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_10_5_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_8_5_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_9_6_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_9_4_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_10_5_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_9_5_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_9_5_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_9_5_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_9_5_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_9_5_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_9_5_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_9_5_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_9_5_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_9_5_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_9_5_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_9_5_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_9_5_out_S_noc3_yummy )
);


tile
tile165 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[165] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd5),
    .default_coreid_y           (8'd10),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd165)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[165]   )
    ,.unavailable_o       ( unavailable_o[165] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[165]   )
    ,.ipi_i               ( ipi_i[165]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[165*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile165_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile165_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_9_5_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_10_6_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_10_4_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_11_5_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_9_5_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_10_6_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_10_4_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_11_5_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_9_5_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_10_6_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_10_4_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_11_5_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_10_5_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_10_5_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_10_5_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_10_5_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_10_5_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_10_5_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_10_5_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_10_5_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_10_5_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_10_5_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_10_5_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_10_5_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_9_5_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_10_6_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_10_4_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_11_5_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_9_5_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_10_6_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_10_4_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_11_5_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_9_5_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_10_6_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_10_4_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_11_5_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_10_5_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_10_5_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_10_5_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_10_5_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_10_5_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_10_5_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_10_5_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_10_5_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_10_5_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_10_5_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_10_5_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_10_5_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_9_5_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_10_6_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_10_4_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_11_5_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_9_5_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_10_6_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_10_4_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_11_5_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_9_5_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_10_6_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_10_4_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_11_5_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_10_5_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_10_5_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_10_5_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_10_5_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_10_5_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_10_5_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_10_5_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_10_5_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_10_5_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_10_5_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_10_5_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_10_5_out_S_noc3_yummy )
);


tile
tile181 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[181] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd5),
    .default_coreid_y           (8'd11),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd181)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[181]   )
    ,.unavailable_o       ( unavailable_o[181] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[181]   )
    ,.ipi_i               ( ipi_i[181]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[181*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile181_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile181_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_10_5_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_11_6_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_11_4_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_12_5_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_10_5_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_11_6_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_11_4_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_12_5_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_10_5_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_11_6_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_11_4_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_12_5_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_11_5_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_11_5_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_11_5_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_11_5_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_11_5_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_11_5_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_11_5_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_11_5_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_11_5_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_11_5_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_11_5_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_11_5_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_10_5_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_11_6_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_11_4_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_12_5_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_10_5_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_11_6_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_11_4_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_12_5_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_10_5_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_11_6_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_11_4_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_12_5_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_11_5_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_11_5_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_11_5_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_11_5_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_11_5_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_11_5_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_11_5_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_11_5_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_11_5_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_11_5_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_11_5_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_11_5_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_10_5_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_11_6_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_11_4_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_12_5_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_10_5_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_11_6_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_11_4_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_12_5_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_10_5_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_11_6_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_11_4_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_12_5_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_11_5_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_11_5_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_11_5_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_11_5_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_11_5_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_11_5_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_11_5_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_11_5_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_11_5_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_11_5_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_11_5_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_11_5_out_S_noc3_yummy )
);


tile
tile197 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[197] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd5),
    .default_coreid_y           (8'd12),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd197)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[197]   )
    ,.unavailable_o       ( unavailable_o[197] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[197]   )
    ,.ipi_i               ( ipi_i[197]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[197*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile197_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile197_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_11_5_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_12_6_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_12_4_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_13_5_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_11_5_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_12_6_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_12_4_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_13_5_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_11_5_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_12_6_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_12_4_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_13_5_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_12_5_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_12_5_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_12_5_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_12_5_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_12_5_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_12_5_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_12_5_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_12_5_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_12_5_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_12_5_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_12_5_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_12_5_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_11_5_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_12_6_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_12_4_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_13_5_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_11_5_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_12_6_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_12_4_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_13_5_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_11_5_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_12_6_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_12_4_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_13_5_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_12_5_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_12_5_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_12_5_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_12_5_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_12_5_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_12_5_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_12_5_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_12_5_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_12_5_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_12_5_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_12_5_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_12_5_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_11_5_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_12_6_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_12_4_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_13_5_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_11_5_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_12_6_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_12_4_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_13_5_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_11_5_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_12_6_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_12_4_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_13_5_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_12_5_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_12_5_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_12_5_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_12_5_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_12_5_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_12_5_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_12_5_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_12_5_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_12_5_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_12_5_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_12_5_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_12_5_out_S_noc3_yummy )
);


tile
tile213 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[213] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd5),
    .default_coreid_y           (8'd13),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd213)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[213]   )
    ,.unavailable_o       ( unavailable_o[213] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[213]   )
    ,.ipi_i               ( ipi_i[213]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[213*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile213_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile213_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_12_5_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_13_6_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_13_4_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_14_5_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_12_5_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_13_6_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_13_4_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_14_5_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_12_5_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_13_6_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_13_4_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_14_5_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_13_5_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_13_5_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_13_5_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_13_5_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_13_5_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_13_5_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_13_5_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_13_5_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_13_5_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_13_5_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_13_5_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_13_5_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_12_5_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_13_6_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_13_4_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_14_5_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_12_5_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_13_6_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_13_4_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_14_5_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_12_5_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_13_6_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_13_4_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_14_5_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_13_5_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_13_5_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_13_5_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_13_5_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_13_5_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_13_5_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_13_5_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_13_5_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_13_5_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_13_5_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_13_5_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_13_5_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_12_5_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_13_6_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_13_4_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_14_5_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_12_5_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_13_6_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_13_4_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_14_5_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_12_5_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_13_6_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_13_4_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_14_5_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_13_5_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_13_5_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_13_5_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_13_5_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_13_5_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_13_5_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_13_5_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_13_5_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_13_5_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_13_5_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_13_5_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_13_5_out_S_noc3_yummy )
);


tile
tile229 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[229] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd5),
    .default_coreid_y           (8'd14),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd229)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[229]   )
    ,.unavailable_o       ( unavailable_o[229] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[229]   )
    ,.ipi_i               ( ipi_i[229]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[229*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile229_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile229_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_13_5_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_14_6_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_14_4_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_15_5_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_13_5_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_14_6_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_14_4_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_15_5_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_13_5_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_14_6_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_14_4_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_15_5_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_14_5_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_14_5_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_14_5_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_14_5_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_14_5_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_14_5_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_14_5_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_14_5_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_14_5_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_14_5_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_14_5_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_14_5_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_13_5_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_14_6_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_14_4_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_15_5_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_13_5_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_14_6_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_14_4_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_15_5_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_13_5_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_14_6_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_14_4_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_15_5_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_14_5_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_14_5_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_14_5_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_14_5_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_14_5_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_14_5_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_14_5_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_14_5_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_14_5_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_14_5_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_14_5_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_14_5_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_13_5_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_14_6_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_14_4_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_15_5_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_13_5_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_14_6_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_14_4_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_15_5_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_13_5_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_14_6_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_14_4_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_15_5_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_14_5_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_14_5_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_14_5_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_14_5_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_14_5_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_14_5_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_14_5_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_14_5_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_14_5_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_14_5_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_14_5_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_14_5_out_S_noc3_yummy )
);


tile
tile245 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[245] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd5),
    .default_coreid_y           (8'd15),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd245)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[245]   )
    ,.unavailable_o       ( unavailable_o[245] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[245]   )
    ,.ipi_i               ( ipi_i[245]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[245*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile245_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile245_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_14_5_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_15_6_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_15_4_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( dummy_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_14_5_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_15_6_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_15_4_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( dummy_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_14_5_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_15_6_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_15_4_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( dummy_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_15_5_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_15_5_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_15_5_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_15_5_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_15_5_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_15_5_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_15_5_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_15_5_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_15_5_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_15_5_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_15_5_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_15_5_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_14_5_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_15_6_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_15_4_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( dummy_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_14_5_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_15_6_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_15_4_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( dummy_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_14_5_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_15_6_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_15_4_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( dummy_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_15_5_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_15_5_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_15_5_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_15_5_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_15_5_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_15_5_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_15_5_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_15_5_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_15_5_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_15_5_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_15_5_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_15_5_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_14_5_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_15_6_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_15_4_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( dummy_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_14_5_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_15_6_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_15_4_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( dummy_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_14_5_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_15_6_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_15_4_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( dummy_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_15_5_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_15_5_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_15_5_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_15_5_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_15_5_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_15_5_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_15_5_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_15_5_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_15_5_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_15_5_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_15_5_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_15_5_out_S_noc3_yummy )
);


tile
tile6 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[6] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd6),
    .default_coreid_y           (8'd0),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd6)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[6]   )
    ,.unavailable_o       ( unavailable_o[6] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[6]   )
    ,.ipi_i               ( ipi_i[6]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[6*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile6_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile6_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( dummy_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_0_7_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_0_5_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_1_6_out_N_noc1_data   ),
    .dyn0_validIn_N      ( dummy_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_0_7_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_0_5_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_1_6_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( dummy_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_0_7_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_0_5_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_1_6_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_0_6_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_0_6_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_0_6_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_0_6_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_0_6_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_0_6_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_0_6_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_0_6_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_0_6_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_0_6_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_0_6_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_0_6_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( dummy_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_0_7_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_0_5_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_1_6_out_N_noc2_data   ),
    .dyn1_validIn_N      ( dummy_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_0_7_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_0_5_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_1_6_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( dummy_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_0_7_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_0_5_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_1_6_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_0_6_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_0_6_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_0_6_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_0_6_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_0_6_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_0_6_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_0_6_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_0_6_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_0_6_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_0_6_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_0_6_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_0_6_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( dummy_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_0_7_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_0_5_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_1_6_out_N_noc3_data   ),
    .dyn2_validIn_N      ( dummy_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_0_7_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_0_5_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_1_6_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( dummy_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_0_7_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_0_5_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_1_6_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_0_6_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_0_6_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_0_6_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_0_6_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_0_6_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_0_6_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_0_6_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_0_6_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_0_6_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_0_6_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_0_6_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_0_6_out_S_noc3_yummy )
);


tile
tile22 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[22] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd6),
    .default_coreid_y           (8'd1),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd22)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[22]   )
    ,.unavailable_o       ( unavailable_o[22] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[22]   )
    ,.ipi_i               ( ipi_i[22]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[22*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile22_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile22_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_0_6_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_1_7_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_1_5_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_2_6_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_0_6_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_1_7_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_1_5_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_2_6_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_0_6_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_1_7_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_1_5_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_2_6_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_1_6_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_1_6_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_1_6_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_1_6_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_1_6_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_1_6_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_1_6_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_1_6_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_1_6_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_1_6_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_1_6_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_1_6_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_0_6_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_1_7_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_1_5_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_2_6_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_0_6_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_1_7_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_1_5_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_2_6_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_0_6_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_1_7_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_1_5_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_2_6_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_1_6_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_1_6_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_1_6_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_1_6_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_1_6_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_1_6_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_1_6_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_1_6_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_1_6_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_1_6_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_1_6_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_1_6_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_0_6_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_1_7_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_1_5_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_2_6_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_0_6_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_1_7_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_1_5_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_2_6_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_0_6_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_1_7_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_1_5_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_2_6_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_1_6_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_1_6_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_1_6_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_1_6_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_1_6_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_1_6_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_1_6_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_1_6_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_1_6_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_1_6_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_1_6_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_1_6_out_S_noc3_yummy )
);


tile
tile38 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[38] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd6),
    .default_coreid_y           (8'd2),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd38)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[38]   )
    ,.unavailable_o       ( unavailable_o[38] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[38]   )
    ,.ipi_i               ( ipi_i[38]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[38*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile38_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile38_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_1_6_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_2_7_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_2_5_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_3_6_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_1_6_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_2_7_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_2_5_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_3_6_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_1_6_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_2_7_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_2_5_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_3_6_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_2_6_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_2_6_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_2_6_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_2_6_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_2_6_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_2_6_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_2_6_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_2_6_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_2_6_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_2_6_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_2_6_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_2_6_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_1_6_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_2_7_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_2_5_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_3_6_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_1_6_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_2_7_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_2_5_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_3_6_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_1_6_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_2_7_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_2_5_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_3_6_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_2_6_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_2_6_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_2_6_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_2_6_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_2_6_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_2_6_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_2_6_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_2_6_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_2_6_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_2_6_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_2_6_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_2_6_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_1_6_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_2_7_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_2_5_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_3_6_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_1_6_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_2_7_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_2_5_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_3_6_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_1_6_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_2_7_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_2_5_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_3_6_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_2_6_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_2_6_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_2_6_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_2_6_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_2_6_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_2_6_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_2_6_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_2_6_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_2_6_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_2_6_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_2_6_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_2_6_out_S_noc3_yummy )
);


tile
tile54 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[54] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd6),
    .default_coreid_y           (8'd3),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd54)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[54]   )
    ,.unavailable_o       ( unavailable_o[54] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[54]   )
    ,.ipi_i               ( ipi_i[54]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[54*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile54_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile54_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_2_6_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_3_7_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_3_5_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_4_6_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_2_6_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_3_7_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_3_5_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_4_6_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_2_6_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_3_7_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_3_5_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_4_6_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_3_6_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_3_6_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_3_6_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_3_6_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_3_6_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_3_6_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_3_6_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_3_6_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_3_6_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_3_6_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_3_6_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_3_6_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_2_6_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_3_7_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_3_5_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_4_6_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_2_6_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_3_7_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_3_5_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_4_6_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_2_6_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_3_7_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_3_5_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_4_6_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_3_6_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_3_6_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_3_6_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_3_6_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_3_6_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_3_6_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_3_6_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_3_6_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_3_6_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_3_6_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_3_6_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_3_6_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_2_6_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_3_7_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_3_5_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_4_6_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_2_6_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_3_7_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_3_5_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_4_6_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_2_6_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_3_7_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_3_5_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_4_6_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_3_6_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_3_6_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_3_6_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_3_6_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_3_6_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_3_6_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_3_6_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_3_6_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_3_6_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_3_6_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_3_6_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_3_6_out_S_noc3_yummy )
);


tile
tile70 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[70] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd6),
    .default_coreid_y           (8'd4),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd70)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[70]   )
    ,.unavailable_o       ( unavailable_o[70] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[70]   )
    ,.ipi_i               ( ipi_i[70]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[70*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile70_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile70_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_3_6_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_4_7_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_4_5_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_5_6_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_3_6_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_4_7_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_4_5_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_5_6_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_3_6_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_4_7_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_4_5_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_5_6_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_4_6_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_4_6_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_4_6_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_4_6_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_4_6_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_4_6_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_4_6_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_4_6_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_4_6_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_4_6_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_4_6_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_4_6_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_3_6_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_4_7_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_4_5_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_5_6_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_3_6_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_4_7_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_4_5_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_5_6_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_3_6_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_4_7_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_4_5_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_5_6_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_4_6_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_4_6_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_4_6_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_4_6_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_4_6_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_4_6_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_4_6_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_4_6_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_4_6_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_4_6_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_4_6_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_4_6_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_3_6_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_4_7_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_4_5_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_5_6_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_3_6_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_4_7_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_4_5_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_5_6_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_3_6_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_4_7_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_4_5_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_5_6_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_4_6_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_4_6_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_4_6_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_4_6_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_4_6_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_4_6_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_4_6_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_4_6_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_4_6_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_4_6_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_4_6_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_4_6_out_S_noc3_yummy )
);


tile
tile86 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[86] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd6),
    .default_coreid_y           (8'd5),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd86)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[86]   )
    ,.unavailable_o       ( unavailable_o[86] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[86]   )
    ,.ipi_i               ( ipi_i[86]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[86*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile86_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile86_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_4_6_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_5_7_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_5_5_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_6_6_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_4_6_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_5_7_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_5_5_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_6_6_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_4_6_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_5_7_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_5_5_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_6_6_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_5_6_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_5_6_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_5_6_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_5_6_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_5_6_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_5_6_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_5_6_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_5_6_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_5_6_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_5_6_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_5_6_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_5_6_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_4_6_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_5_7_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_5_5_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_6_6_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_4_6_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_5_7_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_5_5_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_6_6_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_4_6_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_5_7_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_5_5_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_6_6_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_5_6_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_5_6_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_5_6_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_5_6_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_5_6_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_5_6_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_5_6_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_5_6_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_5_6_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_5_6_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_5_6_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_5_6_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_4_6_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_5_7_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_5_5_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_6_6_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_4_6_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_5_7_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_5_5_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_6_6_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_4_6_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_5_7_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_5_5_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_6_6_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_5_6_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_5_6_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_5_6_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_5_6_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_5_6_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_5_6_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_5_6_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_5_6_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_5_6_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_5_6_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_5_6_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_5_6_out_S_noc3_yummy )
);


tile
tile102 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[102] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd6),
    .default_coreid_y           (8'd6),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd102)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[102]   )
    ,.unavailable_o       ( unavailable_o[102] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[102]   )
    ,.ipi_i               ( ipi_i[102]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[102*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile102_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile102_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_5_6_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_6_7_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_6_5_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_7_6_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_5_6_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_6_7_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_6_5_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_7_6_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_5_6_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_6_7_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_6_5_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_7_6_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_6_6_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_6_6_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_6_6_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_6_6_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_6_6_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_6_6_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_6_6_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_6_6_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_6_6_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_6_6_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_6_6_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_6_6_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_5_6_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_6_7_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_6_5_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_7_6_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_5_6_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_6_7_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_6_5_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_7_6_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_5_6_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_6_7_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_6_5_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_7_6_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_6_6_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_6_6_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_6_6_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_6_6_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_6_6_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_6_6_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_6_6_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_6_6_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_6_6_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_6_6_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_6_6_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_6_6_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_5_6_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_6_7_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_6_5_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_7_6_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_5_6_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_6_7_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_6_5_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_7_6_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_5_6_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_6_7_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_6_5_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_7_6_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_6_6_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_6_6_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_6_6_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_6_6_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_6_6_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_6_6_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_6_6_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_6_6_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_6_6_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_6_6_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_6_6_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_6_6_out_S_noc3_yummy )
);


tile
tile118 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[118] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd6),
    .default_coreid_y           (8'd7),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd118)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[118]   )
    ,.unavailable_o       ( unavailable_o[118] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[118]   )
    ,.ipi_i               ( ipi_i[118]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[118*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile118_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile118_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_6_6_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_7_7_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_7_5_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_8_6_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_6_6_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_7_7_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_7_5_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_8_6_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_6_6_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_7_7_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_7_5_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_8_6_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_7_6_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_7_6_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_7_6_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_7_6_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_7_6_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_7_6_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_7_6_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_7_6_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_7_6_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_7_6_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_7_6_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_7_6_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_6_6_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_7_7_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_7_5_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_8_6_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_6_6_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_7_7_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_7_5_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_8_6_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_6_6_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_7_7_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_7_5_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_8_6_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_7_6_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_7_6_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_7_6_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_7_6_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_7_6_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_7_6_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_7_6_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_7_6_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_7_6_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_7_6_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_7_6_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_7_6_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_6_6_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_7_7_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_7_5_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_8_6_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_6_6_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_7_7_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_7_5_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_8_6_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_6_6_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_7_7_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_7_5_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_8_6_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_7_6_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_7_6_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_7_6_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_7_6_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_7_6_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_7_6_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_7_6_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_7_6_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_7_6_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_7_6_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_7_6_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_7_6_out_S_noc3_yummy )
);


tile
tile134 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[134] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd6),
    .default_coreid_y           (8'd8),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd134)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[134]   )
    ,.unavailable_o       ( unavailable_o[134] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[134]   )
    ,.ipi_i               ( ipi_i[134]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[134*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile134_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile134_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_7_6_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_8_7_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_8_5_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_9_6_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_7_6_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_8_7_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_8_5_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_9_6_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_7_6_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_8_7_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_8_5_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_9_6_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_8_6_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_8_6_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_8_6_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_8_6_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_8_6_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_8_6_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_8_6_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_8_6_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_8_6_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_8_6_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_8_6_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_8_6_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_7_6_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_8_7_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_8_5_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_9_6_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_7_6_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_8_7_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_8_5_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_9_6_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_7_6_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_8_7_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_8_5_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_9_6_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_8_6_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_8_6_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_8_6_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_8_6_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_8_6_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_8_6_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_8_6_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_8_6_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_8_6_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_8_6_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_8_6_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_8_6_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_7_6_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_8_7_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_8_5_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_9_6_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_7_6_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_8_7_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_8_5_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_9_6_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_7_6_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_8_7_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_8_5_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_9_6_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_8_6_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_8_6_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_8_6_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_8_6_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_8_6_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_8_6_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_8_6_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_8_6_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_8_6_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_8_6_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_8_6_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_8_6_out_S_noc3_yummy )
);


tile
tile150 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[150] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd6),
    .default_coreid_y           (8'd9),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd150)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[150]   )
    ,.unavailable_o       ( unavailable_o[150] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[150]   )
    ,.ipi_i               ( ipi_i[150]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[150*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile150_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile150_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_8_6_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_9_7_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_9_5_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_10_6_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_8_6_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_9_7_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_9_5_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_10_6_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_8_6_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_9_7_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_9_5_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_10_6_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_9_6_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_9_6_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_9_6_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_9_6_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_9_6_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_9_6_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_9_6_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_9_6_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_9_6_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_9_6_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_9_6_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_9_6_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_8_6_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_9_7_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_9_5_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_10_6_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_8_6_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_9_7_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_9_5_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_10_6_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_8_6_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_9_7_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_9_5_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_10_6_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_9_6_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_9_6_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_9_6_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_9_6_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_9_6_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_9_6_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_9_6_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_9_6_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_9_6_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_9_6_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_9_6_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_9_6_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_8_6_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_9_7_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_9_5_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_10_6_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_8_6_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_9_7_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_9_5_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_10_6_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_8_6_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_9_7_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_9_5_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_10_6_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_9_6_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_9_6_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_9_6_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_9_6_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_9_6_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_9_6_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_9_6_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_9_6_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_9_6_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_9_6_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_9_6_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_9_6_out_S_noc3_yummy )
);


tile
tile166 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[166] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd6),
    .default_coreid_y           (8'd10),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd166)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[166]   )
    ,.unavailable_o       ( unavailable_o[166] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[166]   )
    ,.ipi_i               ( ipi_i[166]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[166*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile166_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile166_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_9_6_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_10_7_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_10_5_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_11_6_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_9_6_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_10_7_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_10_5_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_11_6_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_9_6_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_10_7_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_10_5_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_11_6_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_10_6_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_10_6_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_10_6_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_10_6_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_10_6_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_10_6_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_10_6_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_10_6_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_10_6_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_10_6_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_10_6_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_10_6_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_9_6_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_10_7_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_10_5_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_11_6_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_9_6_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_10_7_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_10_5_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_11_6_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_9_6_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_10_7_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_10_5_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_11_6_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_10_6_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_10_6_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_10_6_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_10_6_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_10_6_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_10_6_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_10_6_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_10_6_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_10_6_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_10_6_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_10_6_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_10_6_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_9_6_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_10_7_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_10_5_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_11_6_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_9_6_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_10_7_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_10_5_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_11_6_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_9_6_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_10_7_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_10_5_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_11_6_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_10_6_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_10_6_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_10_6_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_10_6_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_10_6_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_10_6_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_10_6_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_10_6_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_10_6_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_10_6_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_10_6_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_10_6_out_S_noc3_yummy )
);


tile
tile182 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[182] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd6),
    .default_coreid_y           (8'd11),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd182)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[182]   )
    ,.unavailable_o       ( unavailable_o[182] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[182]   )
    ,.ipi_i               ( ipi_i[182]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[182*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile182_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile182_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_10_6_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_11_7_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_11_5_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_12_6_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_10_6_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_11_7_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_11_5_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_12_6_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_10_6_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_11_7_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_11_5_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_12_6_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_11_6_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_11_6_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_11_6_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_11_6_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_11_6_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_11_6_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_11_6_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_11_6_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_11_6_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_11_6_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_11_6_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_11_6_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_10_6_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_11_7_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_11_5_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_12_6_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_10_6_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_11_7_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_11_5_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_12_6_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_10_6_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_11_7_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_11_5_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_12_6_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_11_6_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_11_6_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_11_6_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_11_6_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_11_6_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_11_6_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_11_6_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_11_6_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_11_6_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_11_6_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_11_6_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_11_6_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_10_6_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_11_7_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_11_5_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_12_6_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_10_6_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_11_7_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_11_5_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_12_6_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_10_6_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_11_7_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_11_5_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_12_6_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_11_6_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_11_6_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_11_6_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_11_6_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_11_6_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_11_6_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_11_6_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_11_6_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_11_6_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_11_6_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_11_6_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_11_6_out_S_noc3_yummy )
);


tile
tile198 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[198] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd6),
    .default_coreid_y           (8'd12),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd198)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[198]   )
    ,.unavailable_o       ( unavailable_o[198] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[198]   )
    ,.ipi_i               ( ipi_i[198]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[198*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile198_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile198_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_11_6_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_12_7_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_12_5_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_13_6_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_11_6_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_12_7_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_12_5_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_13_6_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_11_6_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_12_7_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_12_5_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_13_6_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_12_6_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_12_6_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_12_6_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_12_6_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_12_6_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_12_6_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_12_6_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_12_6_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_12_6_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_12_6_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_12_6_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_12_6_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_11_6_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_12_7_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_12_5_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_13_6_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_11_6_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_12_7_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_12_5_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_13_6_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_11_6_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_12_7_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_12_5_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_13_6_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_12_6_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_12_6_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_12_6_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_12_6_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_12_6_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_12_6_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_12_6_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_12_6_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_12_6_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_12_6_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_12_6_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_12_6_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_11_6_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_12_7_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_12_5_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_13_6_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_11_6_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_12_7_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_12_5_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_13_6_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_11_6_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_12_7_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_12_5_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_13_6_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_12_6_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_12_6_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_12_6_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_12_6_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_12_6_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_12_6_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_12_6_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_12_6_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_12_6_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_12_6_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_12_6_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_12_6_out_S_noc3_yummy )
);


tile
tile214 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[214] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd6),
    .default_coreid_y           (8'd13),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd214)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[214]   )
    ,.unavailable_o       ( unavailable_o[214] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[214]   )
    ,.ipi_i               ( ipi_i[214]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[214*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile214_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile214_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_12_6_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_13_7_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_13_5_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_14_6_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_12_6_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_13_7_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_13_5_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_14_6_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_12_6_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_13_7_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_13_5_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_14_6_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_13_6_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_13_6_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_13_6_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_13_6_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_13_6_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_13_6_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_13_6_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_13_6_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_13_6_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_13_6_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_13_6_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_13_6_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_12_6_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_13_7_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_13_5_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_14_6_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_12_6_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_13_7_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_13_5_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_14_6_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_12_6_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_13_7_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_13_5_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_14_6_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_13_6_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_13_6_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_13_6_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_13_6_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_13_6_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_13_6_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_13_6_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_13_6_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_13_6_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_13_6_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_13_6_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_13_6_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_12_6_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_13_7_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_13_5_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_14_6_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_12_6_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_13_7_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_13_5_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_14_6_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_12_6_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_13_7_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_13_5_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_14_6_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_13_6_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_13_6_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_13_6_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_13_6_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_13_6_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_13_6_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_13_6_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_13_6_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_13_6_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_13_6_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_13_6_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_13_6_out_S_noc3_yummy )
);


tile
tile230 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[230] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd6),
    .default_coreid_y           (8'd14),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd230)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[230]   )
    ,.unavailable_o       ( unavailable_o[230] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[230]   )
    ,.ipi_i               ( ipi_i[230]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[230*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile230_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile230_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_13_6_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_14_7_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_14_5_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_15_6_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_13_6_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_14_7_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_14_5_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_15_6_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_13_6_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_14_7_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_14_5_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_15_6_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_14_6_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_14_6_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_14_6_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_14_6_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_14_6_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_14_6_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_14_6_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_14_6_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_14_6_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_14_6_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_14_6_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_14_6_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_13_6_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_14_7_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_14_5_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_15_6_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_13_6_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_14_7_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_14_5_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_15_6_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_13_6_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_14_7_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_14_5_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_15_6_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_14_6_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_14_6_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_14_6_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_14_6_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_14_6_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_14_6_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_14_6_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_14_6_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_14_6_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_14_6_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_14_6_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_14_6_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_13_6_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_14_7_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_14_5_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_15_6_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_13_6_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_14_7_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_14_5_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_15_6_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_13_6_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_14_7_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_14_5_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_15_6_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_14_6_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_14_6_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_14_6_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_14_6_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_14_6_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_14_6_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_14_6_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_14_6_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_14_6_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_14_6_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_14_6_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_14_6_out_S_noc3_yummy )
);


tile
tile246 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[246] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd6),
    .default_coreid_y           (8'd15),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd246)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[246]   )
    ,.unavailable_o       ( unavailable_o[246] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[246]   )
    ,.ipi_i               ( ipi_i[246]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[246*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile246_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile246_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_14_6_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_15_7_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_15_5_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( dummy_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_14_6_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_15_7_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_15_5_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( dummy_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_14_6_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_15_7_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_15_5_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( dummy_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_15_6_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_15_6_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_15_6_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_15_6_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_15_6_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_15_6_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_15_6_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_15_6_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_15_6_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_15_6_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_15_6_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_15_6_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_14_6_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_15_7_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_15_5_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( dummy_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_14_6_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_15_7_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_15_5_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( dummy_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_14_6_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_15_7_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_15_5_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( dummy_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_15_6_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_15_6_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_15_6_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_15_6_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_15_6_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_15_6_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_15_6_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_15_6_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_15_6_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_15_6_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_15_6_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_15_6_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_14_6_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_15_7_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_15_5_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( dummy_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_14_6_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_15_7_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_15_5_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( dummy_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_14_6_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_15_7_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_15_5_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( dummy_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_15_6_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_15_6_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_15_6_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_15_6_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_15_6_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_15_6_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_15_6_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_15_6_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_15_6_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_15_6_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_15_6_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_15_6_out_S_noc3_yummy )
);


tile
tile7 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[7] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd7),
    .default_coreid_y           (8'd0),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd7)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[7]   )
    ,.unavailable_o       ( unavailable_o[7] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[7]   )
    ,.ipi_i               ( ipi_i[7]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[7*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile7_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile7_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( dummy_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_0_8_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_0_6_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_1_7_out_N_noc1_data   ),
    .dyn0_validIn_N      ( dummy_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_0_8_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_0_6_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_1_7_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( dummy_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_0_8_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_0_6_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_1_7_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_0_7_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_0_7_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_0_7_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_0_7_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_0_7_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_0_7_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_0_7_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_0_7_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_0_7_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_0_7_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_0_7_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_0_7_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( dummy_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_0_8_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_0_6_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_1_7_out_N_noc2_data   ),
    .dyn1_validIn_N      ( dummy_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_0_8_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_0_6_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_1_7_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( dummy_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_0_8_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_0_6_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_1_7_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_0_7_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_0_7_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_0_7_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_0_7_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_0_7_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_0_7_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_0_7_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_0_7_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_0_7_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_0_7_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_0_7_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_0_7_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( dummy_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_0_8_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_0_6_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_1_7_out_N_noc3_data   ),
    .dyn2_validIn_N      ( dummy_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_0_8_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_0_6_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_1_7_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( dummy_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_0_8_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_0_6_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_1_7_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_0_7_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_0_7_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_0_7_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_0_7_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_0_7_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_0_7_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_0_7_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_0_7_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_0_7_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_0_7_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_0_7_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_0_7_out_S_noc3_yummy )
);


tile
tile23 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[23] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd7),
    .default_coreid_y           (8'd1),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd23)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[23]   )
    ,.unavailable_o       ( unavailable_o[23] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[23]   )
    ,.ipi_i               ( ipi_i[23]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[23*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile23_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile23_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_0_7_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_1_8_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_1_6_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_2_7_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_0_7_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_1_8_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_1_6_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_2_7_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_0_7_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_1_8_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_1_6_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_2_7_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_1_7_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_1_7_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_1_7_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_1_7_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_1_7_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_1_7_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_1_7_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_1_7_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_1_7_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_1_7_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_1_7_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_1_7_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_0_7_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_1_8_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_1_6_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_2_7_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_0_7_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_1_8_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_1_6_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_2_7_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_0_7_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_1_8_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_1_6_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_2_7_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_1_7_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_1_7_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_1_7_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_1_7_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_1_7_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_1_7_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_1_7_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_1_7_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_1_7_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_1_7_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_1_7_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_1_7_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_0_7_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_1_8_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_1_6_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_2_7_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_0_7_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_1_8_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_1_6_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_2_7_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_0_7_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_1_8_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_1_6_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_2_7_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_1_7_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_1_7_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_1_7_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_1_7_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_1_7_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_1_7_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_1_7_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_1_7_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_1_7_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_1_7_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_1_7_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_1_7_out_S_noc3_yummy )
);


tile
tile39 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[39] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd7),
    .default_coreid_y           (8'd2),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd39)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[39]   )
    ,.unavailable_o       ( unavailable_o[39] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[39]   )
    ,.ipi_i               ( ipi_i[39]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[39*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile39_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile39_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_1_7_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_2_8_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_2_6_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_3_7_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_1_7_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_2_8_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_2_6_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_3_7_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_1_7_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_2_8_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_2_6_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_3_7_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_2_7_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_2_7_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_2_7_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_2_7_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_2_7_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_2_7_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_2_7_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_2_7_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_2_7_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_2_7_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_2_7_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_2_7_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_1_7_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_2_8_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_2_6_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_3_7_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_1_7_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_2_8_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_2_6_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_3_7_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_1_7_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_2_8_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_2_6_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_3_7_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_2_7_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_2_7_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_2_7_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_2_7_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_2_7_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_2_7_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_2_7_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_2_7_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_2_7_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_2_7_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_2_7_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_2_7_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_1_7_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_2_8_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_2_6_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_3_7_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_1_7_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_2_8_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_2_6_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_3_7_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_1_7_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_2_8_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_2_6_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_3_7_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_2_7_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_2_7_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_2_7_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_2_7_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_2_7_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_2_7_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_2_7_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_2_7_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_2_7_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_2_7_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_2_7_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_2_7_out_S_noc3_yummy )
);


tile
tile55 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[55] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd7),
    .default_coreid_y           (8'd3),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd55)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[55]   )
    ,.unavailable_o       ( unavailable_o[55] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[55]   )
    ,.ipi_i               ( ipi_i[55]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[55*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile55_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile55_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_2_7_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_3_8_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_3_6_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_4_7_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_2_7_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_3_8_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_3_6_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_4_7_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_2_7_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_3_8_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_3_6_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_4_7_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_3_7_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_3_7_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_3_7_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_3_7_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_3_7_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_3_7_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_3_7_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_3_7_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_3_7_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_3_7_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_3_7_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_3_7_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_2_7_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_3_8_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_3_6_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_4_7_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_2_7_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_3_8_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_3_6_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_4_7_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_2_7_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_3_8_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_3_6_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_4_7_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_3_7_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_3_7_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_3_7_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_3_7_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_3_7_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_3_7_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_3_7_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_3_7_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_3_7_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_3_7_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_3_7_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_3_7_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_2_7_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_3_8_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_3_6_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_4_7_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_2_7_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_3_8_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_3_6_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_4_7_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_2_7_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_3_8_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_3_6_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_4_7_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_3_7_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_3_7_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_3_7_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_3_7_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_3_7_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_3_7_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_3_7_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_3_7_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_3_7_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_3_7_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_3_7_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_3_7_out_S_noc3_yummy )
);


tile
tile71 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[71] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd7),
    .default_coreid_y           (8'd4),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd71)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[71]   )
    ,.unavailable_o       ( unavailable_o[71] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[71]   )
    ,.ipi_i               ( ipi_i[71]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[71*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile71_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile71_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_3_7_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_4_8_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_4_6_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_5_7_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_3_7_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_4_8_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_4_6_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_5_7_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_3_7_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_4_8_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_4_6_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_5_7_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_4_7_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_4_7_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_4_7_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_4_7_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_4_7_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_4_7_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_4_7_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_4_7_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_4_7_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_4_7_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_4_7_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_4_7_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_3_7_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_4_8_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_4_6_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_5_7_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_3_7_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_4_8_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_4_6_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_5_7_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_3_7_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_4_8_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_4_6_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_5_7_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_4_7_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_4_7_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_4_7_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_4_7_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_4_7_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_4_7_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_4_7_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_4_7_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_4_7_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_4_7_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_4_7_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_4_7_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_3_7_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_4_8_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_4_6_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_5_7_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_3_7_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_4_8_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_4_6_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_5_7_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_3_7_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_4_8_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_4_6_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_5_7_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_4_7_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_4_7_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_4_7_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_4_7_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_4_7_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_4_7_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_4_7_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_4_7_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_4_7_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_4_7_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_4_7_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_4_7_out_S_noc3_yummy )
);


tile
tile87 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[87] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd7),
    .default_coreid_y           (8'd5),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd87)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[87]   )
    ,.unavailable_o       ( unavailable_o[87] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[87]   )
    ,.ipi_i               ( ipi_i[87]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[87*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile87_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile87_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_4_7_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_5_8_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_5_6_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_6_7_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_4_7_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_5_8_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_5_6_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_6_7_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_4_7_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_5_8_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_5_6_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_6_7_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_5_7_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_5_7_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_5_7_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_5_7_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_5_7_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_5_7_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_5_7_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_5_7_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_5_7_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_5_7_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_5_7_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_5_7_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_4_7_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_5_8_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_5_6_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_6_7_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_4_7_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_5_8_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_5_6_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_6_7_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_4_7_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_5_8_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_5_6_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_6_7_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_5_7_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_5_7_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_5_7_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_5_7_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_5_7_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_5_7_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_5_7_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_5_7_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_5_7_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_5_7_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_5_7_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_5_7_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_4_7_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_5_8_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_5_6_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_6_7_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_4_7_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_5_8_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_5_6_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_6_7_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_4_7_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_5_8_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_5_6_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_6_7_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_5_7_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_5_7_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_5_7_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_5_7_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_5_7_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_5_7_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_5_7_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_5_7_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_5_7_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_5_7_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_5_7_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_5_7_out_S_noc3_yummy )
);


tile
tile103 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[103] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd7),
    .default_coreid_y           (8'd6),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd103)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[103]   )
    ,.unavailable_o       ( unavailable_o[103] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[103]   )
    ,.ipi_i               ( ipi_i[103]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[103*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile103_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile103_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_5_7_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_6_8_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_6_6_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_7_7_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_5_7_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_6_8_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_6_6_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_7_7_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_5_7_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_6_8_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_6_6_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_7_7_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_6_7_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_6_7_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_6_7_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_6_7_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_6_7_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_6_7_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_6_7_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_6_7_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_6_7_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_6_7_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_6_7_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_6_7_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_5_7_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_6_8_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_6_6_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_7_7_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_5_7_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_6_8_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_6_6_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_7_7_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_5_7_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_6_8_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_6_6_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_7_7_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_6_7_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_6_7_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_6_7_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_6_7_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_6_7_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_6_7_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_6_7_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_6_7_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_6_7_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_6_7_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_6_7_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_6_7_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_5_7_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_6_8_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_6_6_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_7_7_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_5_7_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_6_8_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_6_6_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_7_7_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_5_7_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_6_8_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_6_6_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_7_7_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_6_7_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_6_7_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_6_7_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_6_7_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_6_7_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_6_7_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_6_7_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_6_7_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_6_7_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_6_7_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_6_7_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_6_7_out_S_noc3_yummy )
);


tile
tile119 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[119] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd7),
    .default_coreid_y           (8'd7),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd119)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[119]   )
    ,.unavailable_o       ( unavailable_o[119] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[119]   )
    ,.ipi_i               ( ipi_i[119]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[119*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile119_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile119_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_6_7_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_7_8_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_7_6_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_8_7_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_6_7_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_7_8_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_7_6_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_8_7_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_6_7_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_7_8_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_7_6_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_8_7_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_7_7_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_7_7_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_7_7_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_7_7_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_7_7_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_7_7_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_7_7_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_7_7_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_7_7_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_7_7_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_7_7_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_7_7_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_6_7_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_7_8_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_7_6_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_8_7_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_6_7_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_7_8_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_7_6_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_8_7_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_6_7_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_7_8_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_7_6_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_8_7_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_7_7_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_7_7_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_7_7_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_7_7_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_7_7_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_7_7_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_7_7_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_7_7_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_7_7_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_7_7_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_7_7_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_7_7_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_6_7_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_7_8_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_7_6_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_8_7_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_6_7_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_7_8_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_7_6_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_8_7_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_6_7_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_7_8_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_7_6_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_8_7_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_7_7_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_7_7_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_7_7_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_7_7_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_7_7_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_7_7_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_7_7_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_7_7_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_7_7_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_7_7_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_7_7_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_7_7_out_S_noc3_yummy )
);


tile
tile135 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[135] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd7),
    .default_coreid_y           (8'd8),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd135)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[135]   )
    ,.unavailable_o       ( unavailable_o[135] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[135]   )
    ,.ipi_i               ( ipi_i[135]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[135*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile135_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile135_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_7_7_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_8_8_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_8_6_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_9_7_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_7_7_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_8_8_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_8_6_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_9_7_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_7_7_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_8_8_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_8_6_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_9_7_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_8_7_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_8_7_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_8_7_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_8_7_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_8_7_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_8_7_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_8_7_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_8_7_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_8_7_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_8_7_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_8_7_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_8_7_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_7_7_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_8_8_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_8_6_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_9_7_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_7_7_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_8_8_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_8_6_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_9_7_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_7_7_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_8_8_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_8_6_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_9_7_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_8_7_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_8_7_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_8_7_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_8_7_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_8_7_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_8_7_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_8_7_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_8_7_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_8_7_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_8_7_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_8_7_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_8_7_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_7_7_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_8_8_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_8_6_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_9_7_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_7_7_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_8_8_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_8_6_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_9_7_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_7_7_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_8_8_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_8_6_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_9_7_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_8_7_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_8_7_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_8_7_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_8_7_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_8_7_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_8_7_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_8_7_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_8_7_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_8_7_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_8_7_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_8_7_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_8_7_out_S_noc3_yummy )
);


tile
tile151 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[151] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd7),
    .default_coreid_y           (8'd9),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd151)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[151]   )
    ,.unavailable_o       ( unavailable_o[151] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[151]   )
    ,.ipi_i               ( ipi_i[151]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[151*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile151_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile151_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_8_7_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_9_8_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_9_6_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_10_7_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_8_7_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_9_8_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_9_6_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_10_7_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_8_7_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_9_8_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_9_6_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_10_7_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_9_7_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_9_7_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_9_7_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_9_7_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_9_7_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_9_7_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_9_7_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_9_7_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_9_7_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_9_7_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_9_7_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_9_7_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_8_7_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_9_8_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_9_6_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_10_7_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_8_7_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_9_8_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_9_6_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_10_7_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_8_7_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_9_8_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_9_6_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_10_7_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_9_7_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_9_7_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_9_7_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_9_7_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_9_7_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_9_7_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_9_7_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_9_7_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_9_7_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_9_7_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_9_7_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_9_7_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_8_7_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_9_8_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_9_6_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_10_7_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_8_7_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_9_8_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_9_6_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_10_7_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_8_7_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_9_8_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_9_6_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_10_7_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_9_7_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_9_7_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_9_7_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_9_7_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_9_7_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_9_7_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_9_7_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_9_7_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_9_7_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_9_7_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_9_7_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_9_7_out_S_noc3_yummy )
);


tile
tile167 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[167] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd7),
    .default_coreid_y           (8'd10),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd167)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[167]   )
    ,.unavailable_o       ( unavailable_o[167] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[167]   )
    ,.ipi_i               ( ipi_i[167]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[167*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile167_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile167_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_9_7_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_10_8_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_10_6_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_11_7_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_9_7_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_10_8_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_10_6_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_11_7_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_9_7_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_10_8_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_10_6_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_11_7_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_10_7_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_10_7_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_10_7_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_10_7_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_10_7_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_10_7_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_10_7_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_10_7_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_10_7_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_10_7_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_10_7_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_10_7_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_9_7_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_10_8_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_10_6_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_11_7_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_9_7_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_10_8_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_10_6_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_11_7_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_9_7_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_10_8_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_10_6_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_11_7_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_10_7_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_10_7_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_10_7_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_10_7_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_10_7_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_10_7_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_10_7_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_10_7_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_10_7_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_10_7_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_10_7_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_10_7_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_9_7_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_10_8_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_10_6_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_11_7_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_9_7_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_10_8_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_10_6_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_11_7_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_9_7_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_10_8_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_10_6_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_11_7_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_10_7_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_10_7_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_10_7_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_10_7_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_10_7_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_10_7_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_10_7_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_10_7_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_10_7_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_10_7_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_10_7_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_10_7_out_S_noc3_yummy )
);


tile
tile183 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[183] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd7),
    .default_coreid_y           (8'd11),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd183)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[183]   )
    ,.unavailable_o       ( unavailable_o[183] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[183]   )
    ,.ipi_i               ( ipi_i[183]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[183*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile183_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile183_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_10_7_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_11_8_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_11_6_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_12_7_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_10_7_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_11_8_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_11_6_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_12_7_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_10_7_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_11_8_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_11_6_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_12_7_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_11_7_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_11_7_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_11_7_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_11_7_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_11_7_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_11_7_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_11_7_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_11_7_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_11_7_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_11_7_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_11_7_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_11_7_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_10_7_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_11_8_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_11_6_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_12_7_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_10_7_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_11_8_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_11_6_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_12_7_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_10_7_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_11_8_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_11_6_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_12_7_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_11_7_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_11_7_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_11_7_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_11_7_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_11_7_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_11_7_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_11_7_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_11_7_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_11_7_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_11_7_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_11_7_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_11_7_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_10_7_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_11_8_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_11_6_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_12_7_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_10_7_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_11_8_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_11_6_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_12_7_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_10_7_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_11_8_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_11_6_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_12_7_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_11_7_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_11_7_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_11_7_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_11_7_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_11_7_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_11_7_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_11_7_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_11_7_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_11_7_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_11_7_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_11_7_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_11_7_out_S_noc3_yummy )
);


tile
tile199 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[199] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd7),
    .default_coreid_y           (8'd12),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd199)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[199]   )
    ,.unavailable_o       ( unavailable_o[199] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[199]   )
    ,.ipi_i               ( ipi_i[199]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[199*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile199_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile199_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_11_7_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_12_8_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_12_6_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_13_7_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_11_7_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_12_8_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_12_6_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_13_7_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_11_7_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_12_8_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_12_6_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_13_7_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_12_7_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_12_7_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_12_7_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_12_7_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_12_7_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_12_7_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_12_7_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_12_7_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_12_7_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_12_7_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_12_7_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_12_7_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_11_7_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_12_8_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_12_6_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_13_7_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_11_7_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_12_8_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_12_6_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_13_7_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_11_7_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_12_8_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_12_6_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_13_7_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_12_7_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_12_7_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_12_7_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_12_7_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_12_7_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_12_7_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_12_7_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_12_7_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_12_7_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_12_7_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_12_7_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_12_7_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_11_7_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_12_8_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_12_6_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_13_7_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_11_7_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_12_8_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_12_6_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_13_7_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_11_7_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_12_8_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_12_6_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_13_7_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_12_7_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_12_7_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_12_7_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_12_7_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_12_7_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_12_7_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_12_7_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_12_7_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_12_7_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_12_7_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_12_7_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_12_7_out_S_noc3_yummy )
);


tile
tile215 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[215] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd7),
    .default_coreid_y           (8'd13),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd215)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[215]   )
    ,.unavailable_o       ( unavailable_o[215] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[215]   )
    ,.ipi_i               ( ipi_i[215]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[215*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile215_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile215_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_12_7_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_13_8_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_13_6_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_14_7_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_12_7_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_13_8_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_13_6_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_14_7_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_12_7_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_13_8_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_13_6_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_14_7_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_13_7_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_13_7_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_13_7_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_13_7_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_13_7_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_13_7_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_13_7_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_13_7_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_13_7_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_13_7_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_13_7_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_13_7_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_12_7_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_13_8_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_13_6_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_14_7_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_12_7_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_13_8_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_13_6_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_14_7_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_12_7_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_13_8_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_13_6_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_14_7_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_13_7_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_13_7_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_13_7_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_13_7_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_13_7_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_13_7_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_13_7_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_13_7_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_13_7_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_13_7_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_13_7_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_13_7_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_12_7_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_13_8_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_13_6_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_14_7_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_12_7_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_13_8_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_13_6_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_14_7_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_12_7_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_13_8_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_13_6_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_14_7_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_13_7_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_13_7_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_13_7_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_13_7_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_13_7_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_13_7_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_13_7_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_13_7_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_13_7_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_13_7_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_13_7_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_13_7_out_S_noc3_yummy )
);


tile
tile231 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[231] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd7),
    .default_coreid_y           (8'd14),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd231)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[231]   )
    ,.unavailable_o       ( unavailable_o[231] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[231]   )
    ,.ipi_i               ( ipi_i[231]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[231*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile231_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile231_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_13_7_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_14_8_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_14_6_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_15_7_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_13_7_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_14_8_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_14_6_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_15_7_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_13_7_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_14_8_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_14_6_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_15_7_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_14_7_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_14_7_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_14_7_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_14_7_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_14_7_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_14_7_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_14_7_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_14_7_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_14_7_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_14_7_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_14_7_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_14_7_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_13_7_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_14_8_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_14_6_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_15_7_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_13_7_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_14_8_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_14_6_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_15_7_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_13_7_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_14_8_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_14_6_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_15_7_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_14_7_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_14_7_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_14_7_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_14_7_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_14_7_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_14_7_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_14_7_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_14_7_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_14_7_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_14_7_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_14_7_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_14_7_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_13_7_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_14_8_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_14_6_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_15_7_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_13_7_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_14_8_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_14_6_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_15_7_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_13_7_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_14_8_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_14_6_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_15_7_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_14_7_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_14_7_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_14_7_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_14_7_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_14_7_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_14_7_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_14_7_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_14_7_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_14_7_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_14_7_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_14_7_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_14_7_out_S_noc3_yummy )
);


tile
tile247 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[247] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd7),
    .default_coreid_y           (8'd15),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd247)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[247]   )
    ,.unavailable_o       ( unavailable_o[247] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[247]   )
    ,.ipi_i               ( ipi_i[247]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[247*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile247_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile247_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_14_7_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_15_8_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_15_6_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( dummy_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_14_7_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_15_8_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_15_6_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( dummy_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_14_7_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_15_8_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_15_6_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( dummy_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_15_7_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_15_7_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_15_7_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_15_7_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_15_7_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_15_7_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_15_7_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_15_7_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_15_7_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_15_7_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_15_7_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_15_7_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_14_7_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_15_8_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_15_6_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( dummy_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_14_7_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_15_8_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_15_6_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( dummy_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_14_7_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_15_8_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_15_6_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( dummy_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_15_7_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_15_7_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_15_7_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_15_7_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_15_7_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_15_7_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_15_7_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_15_7_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_15_7_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_15_7_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_15_7_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_15_7_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_14_7_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_15_8_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_15_6_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( dummy_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_14_7_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_15_8_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_15_6_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( dummy_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_14_7_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_15_8_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_15_6_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( dummy_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_15_7_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_15_7_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_15_7_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_15_7_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_15_7_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_15_7_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_15_7_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_15_7_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_15_7_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_15_7_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_15_7_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_15_7_out_S_noc3_yummy )
);


tile
tile8 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[8] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd8),
    .default_coreid_y           (8'd0),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd8)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[8]   )
    ,.unavailable_o       ( unavailable_o[8] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[8]   )
    ,.ipi_i               ( ipi_i[8]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[8*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile8_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile8_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( dummy_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_0_9_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_0_7_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_1_8_out_N_noc1_data   ),
    .dyn0_validIn_N      ( dummy_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_0_9_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_0_7_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_1_8_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( dummy_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_0_9_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_0_7_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_1_8_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_0_8_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_0_8_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_0_8_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_0_8_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_0_8_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_0_8_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_0_8_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_0_8_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_0_8_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_0_8_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_0_8_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_0_8_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( dummy_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_0_9_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_0_7_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_1_8_out_N_noc2_data   ),
    .dyn1_validIn_N      ( dummy_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_0_9_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_0_7_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_1_8_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( dummy_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_0_9_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_0_7_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_1_8_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_0_8_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_0_8_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_0_8_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_0_8_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_0_8_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_0_8_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_0_8_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_0_8_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_0_8_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_0_8_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_0_8_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_0_8_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( dummy_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_0_9_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_0_7_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_1_8_out_N_noc3_data   ),
    .dyn2_validIn_N      ( dummy_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_0_9_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_0_7_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_1_8_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( dummy_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_0_9_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_0_7_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_1_8_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_0_8_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_0_8_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_0_8_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_0_8_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_0_8_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_0_8_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_0_8_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_0_8_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_0_8_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_0_8_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_0_8_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_0_8_out_S_noc3_yummy )
);


tile
tile24 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[24] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd8),
    .default_coreid_y           (8'd1),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd24)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[24]   )
    ,.unavailable_o       ( unavailable_o[24] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[24]   )
    ,.ipi_i               ( ipi_i[24]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[24*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile24_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile24_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_0_8_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_1_9_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_1_7_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_2_8_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_0_8_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_1_9_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_1_7_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_2_8_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_0_8_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_1_9_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_1_7_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_2_8_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_1_8_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_1_8_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_1_8_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_1_8_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_1_8_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_1_8_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_1_8_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_1_8_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_1_8_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_1_8_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_1_8_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_1_8_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_0_8_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_1_9_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_1_7_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_2_8_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_0_8_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_1_9_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_1_7_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_2_8_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_0_8_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_1_9_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_1_7_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_2_8_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_1_8_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_1_8_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_1_8_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_1_8_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_1_8_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_1_8_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_1_8_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_1_8_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_1_8_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_1_8_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_1_8_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_1_8_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_0_8_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_1_9_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_1_7_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_2_8_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_0_8_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_1_9_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_1_7_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_2_8_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_0_8_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_1_9_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_1_7_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_2_8_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_1_8_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_1_8_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_1_8_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_1_8_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_1_8_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_1_8_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_1_8_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_1_8_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_1_8_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_1_8_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_1_8_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_1_8_out_S_noc3_yummy )
);


tile
tile40 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[40] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd8),
    .default_coreid_y           (8'd2),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd40)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[40]   )
    ,.unavailable_o       ( unavailable_o[40] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[40]   )
    ,.ipi_i               ( ipi_i[40]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[40*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile40_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile40_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_1_8_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_2_9_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_2_7_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_3_8_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_1_8_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_2_9_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_2_7_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_3_8_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_1_8_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_2_9_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_2_7_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_3_8_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_2_8_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_2_8_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_2_8_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_2_8_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_2_8_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_2_8_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_2_8_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_2_8_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_2_8_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_2_8_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_2_8_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_2_8_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_1_8_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_2_9_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_2_7_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_3_8_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_1_8_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_2_9_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_2_7_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_3_8_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_1_8_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_2_9_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_2_7_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_3_8_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_2_8_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_2_8_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_2_8_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_2_8_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_2_8_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_2_8_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_2_8_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_2_8_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_2_8_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_2_8_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_2_8_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_2_8_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_1_8_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_2_9_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_2_7_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_3_8_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_1_8_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_2_9_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_2_7_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_3_8_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_1_8_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_2_9_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_2_7_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_3_8_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_2_8_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_2_8_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_2_8_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_2_8_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_2_8_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_2_8_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_2_8_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_2_8_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_2_8_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_2_8_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_2_8_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_2_8_out_S_noc3_yummy )
);


tile
tile56 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[56] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd8),
    .default_coreid_y           (8'd3),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd56)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[56]   )
    ,.unavailable_o       ( unavailable_o[56] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[56]   )
    ,.ipi_i               ( ipi_i[56]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[56*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile56_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile56_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_2_8_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_3_9_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_3_7_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_4_8_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_2_8_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_3_9_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_3_7_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_4_8_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_2_8_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_3_9_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_3_7_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_4_8_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_3_8_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_3_8_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_3_8_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_3_8_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_3_8_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_3_8_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_3_8_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_3_8_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_3_8_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_3_8_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_3_8_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_3_8_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_2_8_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_3_9_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_3_7_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_4_8_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_2_8_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_3_9_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_3_7_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_4_8_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_2_8_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_3_9_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_3_7_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_4_8_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_3_8_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_3_8_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_3_8_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_3_8_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_3_8_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_3_8_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_3_8_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_3_8_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_3_8_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_3_8_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_3_8_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_3_8_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_2_8_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_3_9_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_3_7_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_4_8_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_2_8_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_3_9_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_3_7_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_4_8_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_2_8_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_3_9_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_3_7_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_4_8_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_3_8_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_3_8_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_3_8_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_3_8_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_3_8_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_3_8_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_3_8_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_3_8_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_3_8_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_3_8_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_3_8_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_3_8_out_S_noc3_yummy )
);


tile
tile72 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[72] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd8),
    .default_coreid_y           (8'd4),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd72)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[72]   )
    ,.unavailable_o       ( unavailable_o[72] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[72]   )
    ,.ipi_i               ( ipi_i[72]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[72*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile72_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile72_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_3_8_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_4_9_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_4_7_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_5_8_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_3_8_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_4_9_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_4_7_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_5_8_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_3_8_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_4_9_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_4_7_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_5_8_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_4_8_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_4_8_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_4_8_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_4_8_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_4_8_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_4_8_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_4_8_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_4_8_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_4_8_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_4_8_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_4_8_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_4_8_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_3_8_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_4_9_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_4_7_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_5_8_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_3_8_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_4_9_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_4_7_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_5_8_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_3_8_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_4_9_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_4_7_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_5_8_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_4_8_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_4_8_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_4_8_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_4_8_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_4_8_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_4_8_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_4_8_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_4_8_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_4_8_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_4_8_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_4_8_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_4_8_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_3_8_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_4_9_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_4_7_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_5_8_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_3_8_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_4_9_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_4_7_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_5_8_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_3_8_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_4_9_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_4_7_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_5_8_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_4_8_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_4_8_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_4_8_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_4_8_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_4_8_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_4_8_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_4_8_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_4_8_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_4_8_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_4_8_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_4_8_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_4_8_out_S_noc3_yummy )
);


tile
tile88 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[88] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd8),
    .default_coreid_y           (8'd5),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd88)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[88]   )
    ,.unavailable_o       ( unavailable_o[88] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[88]   )
    ,.ipi_i               ( ipi_i[88]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[88*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile88_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile88_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_4_8_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_5_9_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_5_7_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_6_8_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_4_8_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_5_9_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_5_7_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_6_8_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_4_8_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_5_9_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_5_7_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_6_8_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_5_8_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_5_8_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_5_8_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_5_8_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_5_8_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_5_8_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_5_8_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_5_8_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_5_8_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_5_8_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_5_8_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_5_8_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_4_8_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_5_9_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_5_7_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_6_8_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_4_8_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_5_9_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_5_7_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_6_8_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_4_8_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_5_9_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_5_7_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_6_8_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_5_8_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_5_8_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_5_8_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_5_8_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_5_8_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_5_8_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_5_8_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_5_8_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_5_8_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_5_8_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_5_8_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_5_8_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_4_8_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_5_9_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_5_7_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_6_8_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_4_8_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_5_9_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_5_7_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_6_8_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_4_8_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_5_9_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_5_7_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_6_8_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_5_8_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_5_8_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_5_8_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_5_8_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_5_8_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_5_8_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_5_8_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_5_8_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_5_8_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_5_8_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_5_8_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_5_8_out_S_noc3_yummy )
);


tile
tile104 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[104] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd8),
    .default_coreid_y           (8'd6),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd104)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[104]   )
    ,.unavailable_o       ( unavailable_o[104] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[104]   )
    ,.ipi_i               ( ipi_i[104]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[104*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile104_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile104_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_5_8_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_6_9_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_6_7_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_7_8_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_5_8_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_6_9_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_6_7_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_7_8_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_5_8_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_6_9_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_6_7_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_7_8_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_6_8_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_6_8_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_6_8_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_6_8_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_6_8_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_6_8_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_6_8_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_6_8_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_6_8_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_6_8_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_6_8_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_6_8_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_5_8_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_6_9_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_6_7_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_7_8_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_5_8_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_6_9_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_6_7_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_7_8_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_5_8_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_6_9_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_6_7_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_7_8_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_6_8_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_6_8_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_6_8_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_6_8_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_6_8_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_6_8_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_6_8_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_6_8_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_6_8_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_6_8_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_6_8_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_6_8_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_5_8_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_6_9_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_6_7_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_7_8_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_5_8_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_6_9_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_6_7_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_7_8_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_5_8_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_6_9_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_6_7_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_7_8_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_6_8_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_6_8_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_6_8_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_6_8_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_6_8_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_6_8_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_6_8_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_6_8_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_6_8_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_6_8_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_6_8_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_6_8_out_S_noc3_yummy )
);


tile
tile120 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[120] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd8),
    .default_coreid_y           (8'd7),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd120)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[120]   )
    ,.unavailable_o       ( unavailable_o[120] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[120]   )
    ,.ipi_i               ( ipi_i[120]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[120*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile120_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile120_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_6_8_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_7_9_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_7_7_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_8_8_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_6_8_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_7_9_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_7_7_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_8_8_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_6_8_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_7_9_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_7_7_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_8_8_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_7_8_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_7_8_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_7_8_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_7_8_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_7_8_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_7_8_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_7_8_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_7_8_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_7_8_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_7_8_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_7_8_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_7_8_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_6_8_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_7_9_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_7_7_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_8_8_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_6_8_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_7_9_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_7_7_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_8_8_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_6_8_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_7_9_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_7_7_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_8_8_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_7_8_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_7_8_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_7_8_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_7_8_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_7_8_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_7_8_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_7_8_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_7_8_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_7_8_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_7_8_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_7_8_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_7_8_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_6_8_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_7_9_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_7_7_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_8_8_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_6_8_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_7_9_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_7_7_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_8_8_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_6_8_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_7_9_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_7_7_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_8_8_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_7_8_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_7_8_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_7_8_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_7_8_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_7_8_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_7_8_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_7_8_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_7_8_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_7_8_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_7_8_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_7_8_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_7_8_out_S_noc3_yummy )
);


tile
tile136 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[136] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd8),
    .default_coreid_y           (8'd8),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd136)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[136]   )
    ,.unavailable_o       ( unavailable_o[136] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[136]   )
    ,.ipi_i               ( ipi_i[136]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[136*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile136_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile136_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_7_8_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_8_9_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_8_7_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_9_8_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_7_8_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_8_9_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_8_7_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_9_8_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_7_8_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_8_9_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_8_7_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_9_8_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_8_8_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_8_8_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_8_8_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_8_8_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_8_8_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_8_8_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_8_8_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_8_8_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_8_8_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_8_8_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_8_8_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_8_8_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_7_8_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_8_9_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_8_7_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_9_8_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_7_8_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_8_9_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_8_7_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_9_8_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_7_8_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_8_9_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_8_7_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_9_8_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_8_8_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_8_8_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_8_8_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_8_8_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_8_8_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_8_8_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_8_8_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_8_8_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_8_8_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_8_8_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_8_8_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_8_8_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_7_8_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_8_9_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_8_7_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_9_8_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_7_8_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_8_9_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_8_7_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_9_8_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_7_8_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_8_9_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_8_7_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_9_8_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_8_8_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_8_8_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_8_8_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_8_8_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_8_8_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_8_8_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_8_8_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_8_8_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_8_8_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_8_8_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_8_8_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_8_8_out_S_noc3_yummy )
);


tile
tile152 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[152] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd8),
    .default_coreid_y           (8'd9),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd152)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[152]   )
    ,.unavailable_o       ( unavailable_o[152] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[152]   )
    ,.ipi_i               ( ipi_i[152]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[152*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile152_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile152_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_8_8_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_9_9_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_9_7_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_10_8_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_8_8_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_9_9_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_9_7_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_10_8_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_8_8_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_9_9_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_9_7_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_10_8_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_9_8_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_9_8_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_9_8_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_9_8_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_9_8_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_9_8_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_9_8_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_9_8_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_9_8_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_9_8_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_9_8_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_9_8_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_8_8_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_9_9_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_9_7_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_10_8_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_8_8_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_9_9_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_9_7_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_10_8_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_8_8_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_9_9_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_9_7_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_10_8_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_9_8_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_9_8_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_9_8_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_9_8_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_9_8_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_9_8_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_9_8_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_9_8_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_9_8_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_9_8_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_9_8_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_9_8_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_8_8_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_9_9_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_9_7_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_10_8_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_8_8_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_9_9_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_9_7_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_10_8_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_8_8_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_9_9_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_9_7_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_10_8_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_9_8_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_9_8_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_9_8_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_9_8_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_9_8_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_9_8_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_9_8_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_9_8_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_9_8_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_9_8_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_9_8_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_9_8_out_S_noc3_yummy )
);


tile
tile168 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[168] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd8),
    .default_coreid_y           (8'd10),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd168)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[168]   )
    ,.unavailable_o       ( unavailable_o[168] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[168]   )
    ,.ipi_i               ( ipi_i[168]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[168*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile168_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile168_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_9_8_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_10_9_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_10_7_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_11_8_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_9_8_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_10_9_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_10_7_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_11_8_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_9_8_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_10_9_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_10_7_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_11_8_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_10_8_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_10_8_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_10_8_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_10_8_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_10_8_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_10_8_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_10_8_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_10_8_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_10_8_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_10_8_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_10_8_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_10_8_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_9_8_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_10_9_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_10_7_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_11_8_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_9_8_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_10_9_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_10_7_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_11_8_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_9_8_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_10_9_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_10_7_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_11_8_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_10_8_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_10_8_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_10_8_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_10_8_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_10_8_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_10_8_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_10_8_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_10_8_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_10_8_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_10_8_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_10_8_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_10_8_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_9_8_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_10_9_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_10_7_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_11_8_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_9_8_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_10_9_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_10_7_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_11_8_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_9_8_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_10_9_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_10_7_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_11_8_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_10_8_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_10_8_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_10_8_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_10_8_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_10_8_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_10_8_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_10_8_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_10_8_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_10_8_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_10_8_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_10_8_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_10_8_out_S_noc3_yummy )
);


tile
tile184 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[184] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd8),
    .default_coreid_y           (8'd11),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd184)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[184]   )
    ,.unavailable_o       ( unavailable_o[184] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[184]   )
    ,.ipi_i               ( ipi_i[184]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[184*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile184_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile184_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_10_8_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_11_9_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_11_7_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_12_8_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_10_8_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_11_9_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_11_7_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_12_8_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_10_8_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_11_9_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_11_7_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_12_8_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_11_8_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_11_8_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_11_8_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_11_8_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_11_8_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_11_8_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_11_8_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_11_8_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_11_8_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_11_8_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_11_8_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_11_8_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_10_8_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_11_9_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_11_7_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_12_8_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_10_8_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_11_9_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_11_7_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_12_8_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_10_8_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_11_9_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_11_7_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_12_8_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_11_8_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_11_8_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_11_8_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_11_8_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_11_8_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_11_8_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_11_8_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_11_8_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_11_8_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_11_8_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_11_8_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_11_8_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_10_8_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_11_9_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_11_7_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_12_8_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_10_8_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_11_9_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_11_7_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_12_8_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_10_8_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_11_9_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_11_7_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_12_8_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_11_8_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_11_8_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_11_8_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_11_8_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_11_8_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_11_8_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_11_8_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_11_8_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_11_8_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_11_8_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_11_8_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_11_8_out_S_noc3_yummy )
);


tile
tile200 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[200] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd8),
    .default_coreid_y           (8'd12),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd200)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[200]   )
    ,.unavailable_o       ( unavailable_o[200] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[200]   )
    ,.ipi_i               ( ipi_i[200]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[200*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile200_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile200_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_11_8_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_12_9_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_12_7_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_13_8_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_11_8_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_12_9_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_12_7_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_13_8_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_11_8_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_12_9_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_12_7_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_13_8_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_12_8_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_12_8_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_12_8_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_12_8_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_12_8_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_12_8_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_12_8_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_12_8_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_12_8_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_12_8_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_12_8_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_12_8_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_11_8_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_12_9_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_12_7_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_13_8_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_11_8_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_12_9_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_12_7_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_13_8_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_11_8_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_12_9_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_12_7_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_13_8_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_12_8_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_12_8_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_12_8_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_12_8_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_12_8_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_12_8_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_12_8_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_12_8_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_12_8_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_12_8_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_12_8_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_12_8_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_11_8_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_12_9_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_12_7_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_13_8_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_11_8_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_12_9_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_12_7_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_13_8_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_11_8_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_12_9_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_12_7_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_13_8_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_12_8_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_12_8_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_12_8_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_12_8_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_12_8_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_12_8_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_12_8_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_12_8_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_12_8_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_12_8_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_12_8_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_12_8_out_S_noc3_yummy )
);


tile
tile216 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[216] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd8),
    .default_coreid_y           (8'd13),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd216)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[216]   )
    ,.unavailable_o       ( unavailable_o[216] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[216]   )
    ,.ipi_i               ( ipi_i[216]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[216*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile216_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile216_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_12_8_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_13_9_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_13_7_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_14_8_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_12_8_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_13_9_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_13_7_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_14_8_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_12_8_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_13_9_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_13_7_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_14_8_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_13_8_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_13_8_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_13_8_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_13_8_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_13_8_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_13_8_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_13_8_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_13_8_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_13_8_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_13_8_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_13_8_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_13_8_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_12_8_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_13_9_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_13_7_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_14_8_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_12_8_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_13_9_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_13_7_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_14_8_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_12_8_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_13_9_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_13_7_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_14_8_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_13_8_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_13_8_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_13_8_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_13_8_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_13_8_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_13_8_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_13_8_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_13_8_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_13_8_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_13_8_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_13_8_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_13_8_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_12_8_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_13_9_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_13_7_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_14_8_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_12_8_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_13_9_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_13_7_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_14_8_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_12_8_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_13_9_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_13_7_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_14_8_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_13_8_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_13_8_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_13_8_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_13_8_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_13_8_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_13_8_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_13_8_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_13_8_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_13_8_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_13_8_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_13_8_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_13_8_out_S_noc3_yummy )
);


tile
tile232 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[232] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd8),
    .default_coreid_y           (8'd14),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd232)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[232]   )
    ,.unavailable_o       ( unavailable_o[232] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[232]   )
    ,.ipi_i               ( ipi_i[232]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[232*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile232_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile232_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_13_8_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_14_9_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_14_7_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_15_8_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_13_8_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_14_9_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_14_7_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_15_8_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_13_8_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_14_9_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_14_7_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_15_8_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_14_8_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_14_8_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_14_8_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_14_8_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_14_8_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_14_8_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_14_8_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_14_8_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_14_8_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_14_8_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_14_8_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_14_8_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_13_8_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_14_9_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_14_7_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_15_8_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_13_8_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_14_9_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_14_7_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_15_8_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_13_8_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_14_9_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_14_7_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_15_8_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_14_8_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_14_8_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_14_8_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_14_8_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_14_8_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_14_8_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_14_8_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_14_8_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_14_8_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_14_8_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_14_8_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_14_8_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_13_8_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_14_9_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_14_7_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_15_8_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_13_8_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_14_9_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_14_7_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_15_8_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_13_8_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_14_9_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_14_7_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_15_8_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_14_8_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_14_8_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_14_8_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_14_8_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_14_8_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_14_8_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_14_8_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_14_8_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_14_8_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_14_8_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_14_8_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_14_8_out_S_noc3_yummy )
);


tile
tile248 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[248] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd8),
    .default_coreid_y           (8'd15),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd248)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[248]   )
    ,.unavailable_o       ( unavailable_o[248] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[248]   )
    ,.ipi_i               ( ipi_i[248]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[248*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile248_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile248_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_14_8_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_15_9_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_15_7_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( dummy_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_14_8_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_15_9_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_15_7_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( dummy_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_14_8_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_15_9_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_15_7_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( dummy_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_15_8_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_15_8_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_15_8_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_15_8_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_15_8_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_15_8_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_15_8_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_15_8_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_15_8_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_15_8_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_15_8_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_15_8_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_14_8_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_15_9_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_15_7_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( dummy_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_14_8_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_15_9_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_15_7_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( dummy_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_14_8_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_15_9_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_15_7_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( dummy_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_15_8_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_15_8_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_15_8_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_15_8_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_15_8_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_15_8_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_15_8_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_15_8_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_15_8_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_15_8_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_15_8_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_15_8_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_14_8_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_15_9_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_15_7_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( dummy_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_14_8_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_15_9_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_15_7_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( dummy_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_14_8_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_15_9_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_15_7_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( dummy_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_15_8_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_15_8_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_15_8_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_15_8_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_15_8_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_15_8_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_15_8_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_15_8_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_15_8_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_15_8_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_15_8_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_15_8_out_S_noc3_yummy )
);


tile
tile9 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[9] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd9),
    .default_coreid_y           (8'd0),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd9)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[9]   )
    ,.unavailable_o       ( unavailable_o[9] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[9]   )
    ,.ipi_i               ( ipi_i[9]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[9*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile9_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile9_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( dummy_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_0_10_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_0_8_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_1_9_out_N_noc1_data   ),
    .dyn0_validIn_N      ( dummy_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_0_10_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_0_8_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_1_9_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( dummy_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_0_10_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_0_8_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_1_9_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_0_9_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_0_9_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_0_9_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_0_9_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_0_9_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_0_9_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_0_9_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_0_9_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_0_9_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_0_9_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_0_9_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_0_9_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( dummy_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_0_10_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_0_8_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_1_9_out_N_noc2_data   ),
    .dyn1_validIn_N      ( dummy_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_0_10_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_0_8_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_1_9_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( dummy_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_0_10_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_0_8_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_1_9_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_0_9_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_0_9_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_0_9_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_0_9_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_0_9_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_0_9_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_0_9_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_0_9_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_0_9_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_0_9_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_0_9_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_0_9_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( dummy_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_0_10_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_0_8_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_1_9_out_N_noc3_data   ),
    .dyn2_validIn_N      ( dummy_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_0_10_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_0_8_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_1_9_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( dummy_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_0_10_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_0_8_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_1_9_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_0_9_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_0_9_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_0_9_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_0_9_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_0_9_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_0_9_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_0_9_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_0_9_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_0_9_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_0_9_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_0_9_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_0_9_out_S_noc3_yummy )
);


tile
tile25 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[25] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd9),
    .default_coreid_y           (8'd1),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd25)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[25]   )
    ,.unavailable_o       ( unavailable_o[25] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[25]   )
    ,.ipi_i               ( ipi_i[25]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[25*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile25_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile25_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_0_9_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_1_10_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_1_8_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_2_9_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_0_9_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_1_10_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_1_8_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_2_9_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_0_9_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_1_10_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_1_8_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_2_9_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_1_9_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_1_9_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_1_9_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_1_9_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_1_9_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_1_9_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_1_9_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_1_9_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_1_9_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_1_9_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_1_9_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_1_9_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_0_9_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_1_10_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_1_8_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_2_9_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_0_9_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_1_10_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_1_8_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_2_9_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_0_9_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_1_10_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_1_8_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_2_9_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_1_9_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_1_9_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_1_9_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_1_9_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_1_9_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_1_9_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_1_9_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_1_9_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_1_9_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_1_9_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_1_9_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_1_9_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_0_9_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_1_10_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_1_8_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_2_9_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_0_9_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_1_10_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_1_8_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_2_9_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_0_9_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_1_10_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_1_8_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_2_9_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_1_9_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_1_9_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_1_9_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_1_9_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_1_9_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_1_9_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_1_9_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_1_9_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_1_9_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_1_9_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_1_9_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_1_9_out_S_noc3_yummy )
);


tile
tile41 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[41] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd9),
    .default_coreid_y           (8'd2),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd41)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[41]   )
    ,.unavailable_o       ( unavailable_o[41] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[41]   )
    ,.ipi_i               ( ipi_i[41]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[41*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile41_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile41_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_1_9_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_2_10_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_2_8_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_3_9_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_1_9_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_2_10_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_2_8_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_3_9_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_1_9_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_2_10_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_2_8_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_3_9_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_2_9_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_2_9_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_2_9_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_2_9_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_2_9_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_2_9_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_2_9_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_2_9_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_2_9_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_2_9_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_2_9_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_2_9_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_1_9_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_2_10_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_2_8_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_3_9_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_1_9_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_2_10_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_2_8_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_3_9_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_1_9_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_2_10_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_2_8_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_3_9_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_2_9_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_2_9_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_2_9_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_2_9_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_2_9_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_2_9_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_2_9_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_2_9_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_2_9_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_2_9_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_2_9_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_2_9_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_1_9_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_2_10_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_2_8_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_3_9_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_1_9_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_2_10_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_2_8_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_3_9_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_1_9_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_2_10_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_2_8_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_3_9_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_2_9_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_2_9_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_2_9_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_2_9_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_2_9_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_2_9_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_2_9_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_2_9_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_2_9_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_2_9_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_2_9_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_2_9_out_S_noc3_yummy )
);


tile
tile57 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[57] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd9),
    .default_coreid_y           (8'd3),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd57)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[57]   )
    ,.unavailable_o       ( unavailable_o[57] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[57]   )
    ,.ipi_i               ( ipi_i[57]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[57*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile57_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile57_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_2_9_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_3_10_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_3_8_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_4_9_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_2_9_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_3_10_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_3_8_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_4_9_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_2_9_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_3_10_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_3_8_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_4_9_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_3_9_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_3_9_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_3_9_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_3_9_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_3_9_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_3_9_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_3_9_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_3_9_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_3_9_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_3_9_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_3_9_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_3_9_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_2_9_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_3_10_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_3_8_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_4_9_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_2_9_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_3_10_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_3_8_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_4_9_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_2_9_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_3_10_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_3_8_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_4_9_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_3_9_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_3_9_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_3_9_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_3_9_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_3_9_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_3_9_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_3_9_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_3_9_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_3_9_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_3_9_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_3_9_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_3_9_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_2_9_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_3_10_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_3_8_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_4_9_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_2_9_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_3_10_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_3_8_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_4_9_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_2_9_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_3_10_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_3_8_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_4_9_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_3_9_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_3_9_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_3_9_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_3_9_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_3_9_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_3_9_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_3_9_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_3_9_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_3_9_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_3_9_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_3_9_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_3_9_out_S_noc3_yummy )
);


tile
tile73 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[73] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd9),
    .default_coreid_y           (8'd4),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd73)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[73]   )
    ,.unavailable_o       ( unavailable_o[73] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[73]   )
    ,.ipi_i               ( ipi_i[73]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[73*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile73_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile73_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_3_9_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_4_10_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_4_8_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_5_9_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_3_9_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_4_10_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_4_8_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_5_9_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_3_9_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_4_10_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_4_8_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_5_9_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_4_9_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_4_9_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_4_9_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_4_9_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_4_9_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_4_9_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_4_9_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_4_9_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_4_9_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_4_9_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_4_9_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_4_9_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_3_9_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_4_10_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_4_8_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_5_9_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_3_9_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_4_10_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_4_8_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_5_9_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_3_9_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_4_10_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_4_8_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_5_9_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_4_9_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_4_9_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_4_9_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_4_9_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_4_9_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_4_9_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_4_9_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_4_9_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_4_9_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_4_9_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_4_9_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_4_9_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_3_9_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_4_10_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_4_8_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_5_9_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_3_9_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_4_10_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_4_8_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_5_9_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_3_9_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_4_10_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_4_8_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_5_9_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_4_9_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_4_9_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_4_9_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_4_9_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_4_9_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_4_9_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_4_9_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_4_9_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_4_9_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_4_9_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_4_9_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_4_9_out_S_noc3_yummy )
);


tile
tile89 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[89] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd9),
    .default_coreid_y           (8'd5),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd89)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[89]   )
    ,.unavailable_o       ( unavailable_o[89] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[89]   )
    ,.ipi_i               ( ipi_i[89]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[89*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile89_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile89_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_4_9_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_5_10_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_5_8_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_6_9_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_4_9_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_5_10_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_5_8_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_6_9_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_4_9_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_5_10_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_5_8_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_6_9_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_5_9_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_5_9_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_5_9_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_5_9_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_5_9_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_5_9_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_5_9_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_5_9_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_5_9_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_5_9_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_5_9_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_5_9_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_4_9_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_5_10_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_5_8_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_6_9_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_4_9_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_5_10_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_5_8_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_6_9_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_4_9_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_5_10_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_5_8_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_6_9_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_5_9_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_5_9_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_5_9_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_5_9_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_5_9_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_5_9_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_5_9_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_5_9_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_5_9_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_5_9_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_5_9_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_5_9_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_4_9_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_5_10_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_5_8_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_6_9_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_4_9_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_5_10_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_5_8_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_6_9_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_4_9_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_5_10_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_5_8_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_6_9_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_5_9_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_5_9_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_5_9_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_5_9_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_5_9_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_5_9_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_5_9_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_5_9_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_5_9_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_5_9_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_5_9_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_5_9_out_S_noc3_yummy )
);


tile
tile105 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[105] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd9),
    .default_coreid_y           (8'd6),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd105)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[105]   )
    ,.unavailable_o       ( unavailable_o[105] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[105]   )
    ,.ipi_i               ( ipi_i[105]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[105*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile105_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile105_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_5_9_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_6_10_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_6_8_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_7_9_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_5_9_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_6_10_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_6_8_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_7_9_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_5_9_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_6_10_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_6_8_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_7_9_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_6_9_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_6_9_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_6_9_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_6_9_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_6_9_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_6_9_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_6_9_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_6_9_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_6_9_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_6_9_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_6_9_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_6_9_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_5_9_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_6_10_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_6_8_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_7_9_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_5_9_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_6_10_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_6_8_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_7_9_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_5_9_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_6_10_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_6_8_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_7_9_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_6_9_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_6_9_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_6_9_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_6_9_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_6_9_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_6_9_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_6_9_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_6_9_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_6_9_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_6_9_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_6_9_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_6_9_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_5_9_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_6_10_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_6_8_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_7_9_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_5_9_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_6_10_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_6_8_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_7_9_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_5_9_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_6_10_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_6_8_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_7_9_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_6_9_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_6_9_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_6_9_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_6_9_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_6_9_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_6_9_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_6_9_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_6_9_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_6_9_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_6_9_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_6_9_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_6_9_out_S_noc3_yummy )
);


tile
tile121 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[121] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd9),
    .default_coreid_y           (8'd7),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd121)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[121]   )
    ,.unavailable_o       ( unavailable_o[121] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[121]   )
    ,.ipi_i               ( ipi_i[121]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[121*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile121_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile121_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_6_9_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_7_10_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_7_8_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_8_9_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_6_9_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_7_10_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_7_8_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_8_9_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_6_9_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_7_10_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_7_8_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_8_9_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_7_9_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_7_9_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_7_9_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_7_9_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_7_9_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_7_9_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_7_9_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_7_9_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_7_9_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_7_9_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_7_9_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_7_9_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_6_9_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_7_10_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_7_8_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_8_9_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_6_9_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_7_10_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_7_8_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_8_9_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_6_9_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_7_10_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_7_8_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_8_9_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_7_9_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_7_9_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_7_9_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_7_9_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_7_9_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_7_9_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_7_9_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_7_9_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_7_9_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_7_9_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_7_9_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_7_9_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_6_9_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_7_10_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_7_8_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_8_9_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_6_9_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_7_10_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_7_8_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_8_9_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_6_9_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_7_10_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_7_8_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_8_9_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_7_9_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_7_9_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_7_9_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_7_9_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_7_9_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_7_9_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_7_9_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_7_9_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_7_9_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_7_9_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_7_9_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_7_9_out_S_noc3_yummy )
);


tile
tile137 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[137] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd9),
    .default_coreid_y           (8'd8),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd137)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[137]   )
    ,.unavailable_o       ( unavailable_o[137] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[137]   )
    ,.ipi_i               ( ipi_i[137]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[137*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile137_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile137_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_7_9_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_8_10_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_8_8_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_9_9_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_7_9_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_8_10_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_8_8_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_9_9_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_7_9_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_8_10_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_8_8_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_9_9_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_8_9_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_8_9_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_8_9_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_8_9_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_8_9_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_8_9_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_8_9_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_8_9_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_8_9_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_8_9_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_8_9_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_8_9_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_7_9_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_8_10_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_8_8_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_9_9_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_7_9_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_8_10_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_8_8_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_9_9_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_7_9_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_8_10_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_8_8_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_9_9_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_8_9_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_8_9_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_8_9_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_8_9_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_8_9_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_8_9_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_8_9_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_8_9_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_8_9_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_8_9_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_8_9_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_8_9_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_7_9_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_8_10_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_8_8_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_9_9_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_7_9_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_8_10_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_8_8_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_9_9_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_7_9_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_8_10_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_8_8_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_9_9_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_8_9_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_8_9_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_8_9_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_8_9_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_8_9_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_8_9_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_8_9_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_8_9_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_8_9_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_8_9_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_8_9_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_8_9_out_S_noc3_yummy )
);


tile
tile153 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[153] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd9),
    .default_coreid_y           (8'd9),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd153)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[153]   )
    ,.unavailable_o       ( unavailable_o[153] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[153]   )
    ,.ipi_i               ( ipi_i[153]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[153*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile153_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile153_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_8_9_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_9_10_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_9_8_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_10_9_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_8_9_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_9_10_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_9_8_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_10_9_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_8_9_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_9_10_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_9_8_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_10_9_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_9_9_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_9_9_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_9_9_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_9_9_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_9_9_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_9_9_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_9_9_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_9_9_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_9_9_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_9_9_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_9_9_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_9_9_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_8_9_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_9_10_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_9_8_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_10_9_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_8_9_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_9_10_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_9_8_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_10_9_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_8_9_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_9_10_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_9_8_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_10_9_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_9_9_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_9_9_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_9_9_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_9_9_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_9_9_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_9_9_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_9_9_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_9_9_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_9_9_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_9_9_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_9_9_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_9_9_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_8_9_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_9_10_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_9_8_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_10_9_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_8_9_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_9_10_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_9_8_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_10_9_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_8_9_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_9_10_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_9_8_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_10_9_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_9_9_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_9_9_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_9_9_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_9_9_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_9_9_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_9_9_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_9_9_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_9_9_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_9_9_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_9_9_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_9_9_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_9_9_out_S_noc3_yummy )
);


tile
tile169 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[169] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd9),
    .default_coreid_y           (8'd10),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd169)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[169]   )
    ,.unavailable_o       ( unavailable_o[169] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[169]   )
    ,.ipi_i               ( ipi_i[169]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[169*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile169_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile169_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_9_9_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_10_10_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_10_8_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_11_9_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_9_9_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_10_10_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_10_8_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_11_9_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_9_9_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_10_10_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_10_8_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_11_9_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_10_9_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_10_9_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_10_9_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_10_9_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_10_9_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_10_9_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_10_9_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_10_9_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_10_9_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_10_9_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_10_9_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_10_9_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_9_9_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_10_10_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_10_8_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_11_9_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_9_9_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_10_10_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_10_8_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_11_9_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_9_9_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_10_10_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_10_8_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_11_9_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_10_9_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_10_9_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_10_9_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_10_9_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_10_9_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_10_9_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_10_9_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_10_9_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_10_9_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_10_9_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_10_9_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_10_9_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_9_9_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_10_10_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_10_8_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_11_9_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_9_9_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_10_10_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_10_8_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_11_9_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_9_9_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_10_10_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_10_8_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_11_9_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_10_9_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_10_9_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_10_9_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_10_9_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_10_9_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_10_9_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_10_9_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_10_9_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_10_9_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_10_9_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_10_9_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_10_9_out_S_noc3_yummy )
);


tile
tile185 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[185] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd9),
    .default_coreid_y           (8'd11),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd185)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[185]   )
    ,.unavailable_o       ( unavailable_o[185] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[185]   )
    ,.ipi_i               ( ipi_i[185]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[185*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile185_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile185_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_10_9_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_11_10_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_11_8_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_12_9_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_10_9_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_11_10_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_11_8_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_12_9_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_10_9_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_11_10_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_11_8_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_12_9_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_11_9_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_11_9_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_11_9_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_11_9_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_11_9_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_11_9_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_11_9_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_11_9_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_11_9_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_11_9_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_11_9_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_11_9_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_10_9_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_11_10_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_11_8_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_12_9_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_10_9_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_11_10_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_11_8_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_12_9_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_10_9_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_11_10_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_11_8_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_12_9_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_11_9_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_11_9_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_11_9_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_11_9_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_11_9_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_11_9_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_11_9_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_11_9_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_11_9_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_11_9_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_11_9_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_11_9_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_10_9_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_11_10_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_11_8_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_12_9_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_10_9_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_11_10_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_11_8_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_12_9_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_10_9_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_11_10_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_11_8_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_12_9_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_11_9_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_11_9_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_11_9_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_11_9_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_11_9_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_11_9_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_11_9_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_11_9_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_11_9_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_11_9_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_11_9_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_11_9_out_S_noc3_yummy )
);


tile
tile201 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[201] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd9),
    .default_coreid_y           (8'd12),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd201)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[201]   )
    ,.unavailable_o       ( unavailable_o[201] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[201]   )
    ,.ipi_i               ( ipi_i[201]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[201*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile201_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile201_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_11_9_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_12_10_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_12_8_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_13_9_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_11_9_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_12_10_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_12_8_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_13_9_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_11_9_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_12_10_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_12_8_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_13_9_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_12_9_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_12_9_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_12_9_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_12_9_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_12_9_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_12_9_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_12_9_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_12_9_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_12_9_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_12_9_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_12_9_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_12_9_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_11_9_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_12_10_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_12_8_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_13_9_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_11_9_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_12_10_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_12_8_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_13_9_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_11_9_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_12_10_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_12_8_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_13_9_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_12_9_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_12_9_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_12_9_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_12_9_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_12_9_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_12_9_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_12_9_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_12_9_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_12_9_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_12_9_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_12_9_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_12_9_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_11_9_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_12_10_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_12_8_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_13_9_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_11_9_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_12_10_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_12_8_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_13_9_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_11_9_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_12_10_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_12_8_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_13_9_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_12_9_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_12_9_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_12_9_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_12_9_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_12_9_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_12_9_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_12_9_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_12_9_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_12_9_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_12_9_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_12_9_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_12_9_out_S_noc3_yummy )
);


tile
tile217 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[217] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd9),
    .default_coreid_y           (8'd13),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd217)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[217]   )
    ,.unavailable_o       ( unavailable_o[217] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[217]   )
    ,.ipi_i               ( ipi_i[217]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[217*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile217_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile217_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_12_9_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_13_10_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_13_8_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_14_9_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_12_9_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_13_10_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_13_8_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_14_9_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_12_9_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_13_10_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_13_8_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_14_9_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_13_9_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_13_9_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_13_9_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_13_9_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_13_9_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_13_9_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_13_9_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_13_9_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_13_9_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_13_9_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_13_9_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_13_9_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_12_9_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_13_10_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_13_8_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_14_9_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_12_9_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_13_10_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_13_8_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_14_9_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_12_9_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_13_10_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_13_8_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_14_9_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_13_9_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_13_9_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_13_9_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_13_9_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_13_9_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_13_9_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_13_9_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_13_9_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_13_9_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_13_9_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_13_9_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_13_9_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_12_9_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_13_10_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_13_8_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_14_9_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_12_9_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_13_10_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_13_8_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_14_9_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_12_9_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_13_10_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_13_8_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_14_9_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_13_9_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_13_9_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_13_9_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_13_9_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_13_9_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_13_9_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_13_9_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_13_9_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_13_9_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_13_9_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_13_9_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_13_9_out_S_noc3_yummy )
);


tile
tile233 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[233] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd9),
    .default_coreid_y           (8'd14),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd233)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[233]   )
    ,.unavailable_o       ( unavailable_o[233] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[233]   )
    ,.ipi_i               ( ipi_i[233]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[233*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile233_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile233_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_13_9_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_14_10_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_14_8_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_15_9_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_13_9_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_14_10_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_14_8_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_15_9_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_13_9_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_14_10_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_14_8_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_15_9_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_14_9_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_14_9_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_14_9_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_14_9_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_14_9_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_14_9_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_14_9_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_14_9_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_14_9_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_14_9_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_14_9_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_14_9_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_13_9_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_14_10_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_14_8_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_15_9_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_13_9_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_14_10_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_14_8_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_15_9_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_13_9_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_14_10_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_14_8_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_15_9_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_14_9_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_14_9_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_14_9_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_14_9_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_14_9_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_14_9_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_14_9_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_14_9_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_14_9_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_14_9_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_14_9_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_14_9_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_13_9_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_14_10_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_14_8_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_15_9_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_13_9_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_14_10_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_14_8_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_15_9_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_13_9_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_14_10_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_14_8_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_15_9_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_14_9_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_14_9_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_14_9_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_14_9_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_14_9_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_14_9_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_14_9_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_14_9_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_14_9_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_14_9_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_14_9_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_14_9_out_S_noc3_yummy )
);


tile
tile249 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[249] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd9),
    .default_coreid_y           (8'd15),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd249)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[249]   )
    ,.unavailable_o       ( unavailable_o[249] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[249]   )
    ,.ipi_i               ( ipi_i[249]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[249*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile249_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile249_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_14_9_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_15_10_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_15_8_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( dummy_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_14_9_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_15_10_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_15_8_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( dummy_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_14_9_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_15_10_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_15_8_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( dummy_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_15_9_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_15_9_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_15_9_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_15_9_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_15_9_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_15_9_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_15_9_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_15_9_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_15_9_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_15_9_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_15_9_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_15_9_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_14_9_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_15_10_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_15_8_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( dummy_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_14_9_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_15_10_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_15_8_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( dummy_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_14_9_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_15_10_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_15_8_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( dummy_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_15_9_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_15_9_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_15_9_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_15_9_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_15_9_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_15_9_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_15_9_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_15_9_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_15_9_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_15_9_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_15_9_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_15_9_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_14_9_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_15_10_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_15_8_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( dummy_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_14_9_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_15_10_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_15_8_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( dummy_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_14_9_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_15_10_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_15_8_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( dummy_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_15_9_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_15_9_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_15_9_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_15_9_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_15_9_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_15_9_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_15_9_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_15_9_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_15_9_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_15_9_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_15_9_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_15_9_out_S_noc3_yummy )
);


tile
tile10 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[10] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd10),
    .default_coreid_y           (8'd0),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd10)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[10]   )
    ,.unavailable_o       ( unavailable_o[10] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[10]   )
    ,.ipi_i               ( ipi_i[10]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[10*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile10_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile10_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( dummy_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_0_11_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_0_9_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_1_10_out_N_noc1_data   ),
    .dyn0_validIn_N      ( dummy_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_0_11_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_0_9_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_1_10_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( dummy_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_0_11_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_0_9_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_1_10_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_0_10_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_0_10_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_0_10_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_0_10_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_0_10_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_0_10_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_0_10_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_0_10_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_0_10_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_0_10_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_0_10_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_0_10_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( dummy_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_0_11_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_0_9_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_1_10_out_N_noc2_data   ),
    .dyn1_validIn_N      ( dummy_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_0_11_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_0_9_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_1_10_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( dummy_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_0_11_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_0_9_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_1_10_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_0_10_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_0_10_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_0_10_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_0_10_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_0_10_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_0_10_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_0_10_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_0_10_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_0_10_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_0_10_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_0_10_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_0_10_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( dummy_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_0_11_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_0_9_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_1_10_out_N_noc3_data   ),
    .dyn2_validIn_N      ( dummy_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_0_11_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_0_9_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_1_10_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( dummy_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_0_11_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_0_9_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_1_10_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_0_10_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_0_10_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_0_10_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_0_10_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_0_10_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_0_10_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_0_10_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_0_10_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_0_10_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_0_10_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_0_10_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_0_10_out_S_noc3_yummy )
);


tile
tile26 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[26] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd10),
    .default_coreid_y           (8'd1),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd26)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[26]   )
    ,.unavailable_o       ( unavailable_o[26] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[26]   )
    ,.ipi_i               ( ipi_i[26]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[26*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile26_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile26_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_0_10_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_1_11_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_1_9_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_2_10_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_0_10_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_1_11_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_1_9_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_2_10_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_0_10_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_1_11_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_1_9_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_2_10_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_1_10_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_1_10_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_1_10_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_1_10_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_1_10_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_1_10_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_1_10_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_1_10_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_1_10_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_1_10_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_1_10_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_1_10_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_0_10_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_1_11_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_1_9_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_2_10_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_0_10_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_1_11_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_1_9_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_2_10_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_0_10_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_1_11_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_1_9_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_2_10_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_1_10_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_1_10_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_1_10_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_1_10_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_1_10_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_1_10_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_1_10_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_1_10_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_1_10_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_1_10_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_1_10_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_1_10_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_0_10_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_1_11_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_1_9_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_2_10_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_0_10_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_1_11_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_1_9_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_2_10_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_0_10_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_1_11_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_1_9_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_2_10_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_1_10_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_1_10_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_1_10_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_1_10_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_1_10_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_1_10_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_1_10_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_1_10_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_1_10_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_1_10_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_1_10_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_1_10_out_S_noc3_yummy )
);


tile
tile42 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[42] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd10),
    .default_coreid_y           (8'd2),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd42)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[42]   )
    ,.unavailable_o       ( unavailable_o[42] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[42]   )
    ,.ipi_i               ( ipi_i[42]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[42*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile42_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile42_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_1_10_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_2_11_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_2_9_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_3_10_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_1_10_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_2_11_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_2_9_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_3_10_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_1_10_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_2_11_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_2_9_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_3_10_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_2_10_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_2_10_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_2_10_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_2_10_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_2_10_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_2_10_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_2_10_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_2_10_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_2_10_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_2_10_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_2_10_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_2_10_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_1_10_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_2_11_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_2_9_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_3_10_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_1_10_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_2_11_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_2_9_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_3_10_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_1_10_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_2_11_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_2_9_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_3_10_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_2_10_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_2_10_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_2_10_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_2_10_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_2_10_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_2_10_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_2_10_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_2_10_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_2_10_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_2_10_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_2_10_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_2_10_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_1_10_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_2_11_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_2_9_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_3_10_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_1_10_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_2_11_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_2_9_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_3_10_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_1_10_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_2_11_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_2_9_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_3_10_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_2_10_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_2_10_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_2_10_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_2_10_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_2_10_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_2_10_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_2_10_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_2_10_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_2_10_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_2_10_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_2_10_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_2_10_out_S_noc3_yummy )
);


tile
tile58 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[58] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd10),
    .default_coreid_y           (8'd3),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd58)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[58]   )
    ,.unavailable_o       ( unavailable_o[58] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[58]   )
    ,.ipi_i               ( ipi_i[58]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[58*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile58_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile58_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_2_10_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_3_11_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_3_9_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_4_10_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_2_10_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_3_11_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_3_9_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_4_10_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_2_10_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_3_11_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_3_9_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_4_10_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_3_10_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_3_10_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_3_10_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_3_10_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_3_10_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_3_10_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_3_10_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_3_10_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_3_10_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_3_10_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_3_10_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_3_10_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_2_10_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_3_11_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_3_9_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_4_10_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_2_10_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_3_11_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_3_9_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_4_10_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_2_10_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_3_11_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_3_9_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_4_10_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_3_10_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_3_10_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_3_10_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_3_10_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_3_10_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_3_10_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_3_10_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_3_10_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_3_10_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_3_10_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_3_10_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_3_10_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_2_10_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_3_11_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_3_9_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_4_10_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_2_10_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_3_11_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_3_9_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_4_10_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_2_10_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_3_11_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_3_9_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_4_10_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_3_10_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_3_10_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_3_10_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_3_10_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_3_10_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_3_10_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_3_10_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_3_10_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_3_10_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_3_10_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_3_10_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_3_10_out_S_noc3_yummy )
);


tile
tile74 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[74] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd10),
    .default_coreid_y           (8'd4),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd74)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[74]   )
    ,.unavailable_o       ( unavailable_o[74] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[74]   )
    ,.ipi_i               ( ipi_i[74]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[74*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile74_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile74_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_3_10_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_4_11_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_4_9_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_5_10_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_3_10_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_4_11_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_4_9_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_5_10_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_3_10_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_4_11_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_4_9_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_5_10_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_4_10_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_4_10_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_4_10_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_4_10_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_4_10_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_4_10_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_4_10_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_4_10_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_4_10_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_4_10_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_4_10_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_4_10_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_3_10_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_4_11_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_4_9_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_5_10_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_3_10_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_4_11_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_4_9_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_5_10_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_3_10_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_4_11_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_4_9_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_5_10_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_4_10_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_4_10_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_4_10_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_4_10_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_4_10_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_4_10_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_4_10_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_4_10_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_4_10_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_4_10_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_4_10_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_4_10_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_3_10_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_4_11_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_4_9_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_5_10_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_3_10_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_4_11_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_4_9_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_5_10_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_3_10_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_4_11_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_4_9_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_5_10_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_4_10_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_4_10_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_4_10_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_4_10_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_4_10_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_4_10_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_4_10_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_4_10_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_4_10_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_4_10_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_4_10_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_4_10_out_S_noc3_yummy )
);


tile
tile90 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[90] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd10),
    .default_coreid_y           (8'd5),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd90)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[90]   )
    ,.unavailable_o       ( unavailable_o[90] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[90]   )
    ,.ipi_i               ( ipi_i[90]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[90*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile90_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile90_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_4_10_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_5_11_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_5_9_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_6_10_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_4_10_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_5_11_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_5_9_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_6_10_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_4_10_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_5_11_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_5_9_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_6_10_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_5_10_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_5_10_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_5_10_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_5_10_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_5_10_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_5_10_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_5_10_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_5_10_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_5_10_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_5_10_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_5_10_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_5_10_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_4_10_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_5_11_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_5_9_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_6_10_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_4_10_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_5_11_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_5_9_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_6_10_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_4_10_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_5_11_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_5_9_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_6_10_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_5_10_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_5_10_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_5_10_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_5_10_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_5_10_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_5_10_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_5_10_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_5_10_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_5_10_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_5_10_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_5_10_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_5_10_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_4_10_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_5_11_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_5_9_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_6_10_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_4_10_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_5_11_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_5_9_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_6_10_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_4_10_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_5_11_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_5_9_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_6_10_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_5_10_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_5_10_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_5_10_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_5_10_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_5_10_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_5_10_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_5_10_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_5_10_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_5_10_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_5_10_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_5_10_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_5_10_out_S_noc3_yummy )
);


tile
tile106 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[106] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd10),
    .default_coreid_y           (8'd6),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd106)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[106]   )
    ,.unavailable_o       ( unavailable_o[106] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[106]   )
    ,.ipi_i               ( ipi_i[106]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[106*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile106_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile106_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_5_10_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_6_11_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_6_9_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_7_10_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_5_10_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_6_11_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_6_9_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_7_10_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_5_10_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_6_11_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_6_9_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_7_10_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_6_10_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_6_10_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_6_10_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_6_10_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_6_10_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_6_10_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_6_10_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_6_10_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_6_10_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_6_10_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_6_10_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_6_10_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_5_10_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_6_11_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_6_9_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_7_10_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_5_10_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_6_11_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_6_9_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_7_10_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_5_10_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_6_11_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_6_9_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_7_10_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_6_10_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_6_10_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_6_10_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_6_10_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_6_10_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_6_10_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_6_10_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_6_10_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_6_10_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_6_10_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_6_10_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_6_10_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_5_10_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_6_11_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_6_9_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_7_10_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_5_10_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_6_11_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_6_9_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_7_10_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_5_10_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_6_11_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_6_9_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_7_10_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_6_10_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_6_10_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_6_10_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_6_10_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_6_10_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_6_10_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_6_10_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_6_10_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_6_10_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_6_10_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_6_10_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_6_10_out_S_noc3_yummy )
);


tile
tile122 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[122] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd10),
    .default_coreid_y           (8'd7),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd122)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[122]   )
    ,.unavailable_o       ( unavailable_o[122] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[122]   )
    ,.ipi_i               ( ipi_i[122]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[122*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile122_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile122_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_6_10_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_7_11_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_7_9_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_8_10_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_6_10_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_7_11_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_7_9_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_8_10_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_6_10_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_7_11_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_7_9_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_8_10_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_7_10_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_7_10_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_7_10_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_7_10_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_7_10_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_7_10_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_7_10_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_7_10_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_7_10_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_7_10_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_7_10_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_7_10_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_6_10_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_7_11_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_7_9_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_8_10_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_6_10_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_7_11_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_7_9_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_8_10_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_6_10_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_7_11_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_7_9_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_8_10_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_7_10_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_7_10_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_7_10_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_7_10_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_7_10_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_7_10_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_7_10_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_7_10_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_7_10_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_7_10_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_7_10_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_7_10_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_6_10_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_7_11_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_7_9_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_8_10_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_6_10_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_7_11_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_7_9_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_8_10_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_6_10_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_7_11_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_7_9_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_8_10_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_7_10_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_7_10_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_7_10_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_7_10_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_7_10_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_7_10_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_7_10_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_7_10_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_7_10_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_7_10_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_7_10_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_7_10_out_S_noc3_yummy )
);


tile
tile138 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[138] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd10),
    .default_coreid_y           (8'd8),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd138)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[138]   )
    ,.unavailable_o       ( unavailable_o[138] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[138]   )
    ,.ipi_i               ( ipi_i[138]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[138*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile138_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile138_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_7_10_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_8_11_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_8_9_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_9_10_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_7_10_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_8_11_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_8_9_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_9_10_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_7_10_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_8_11_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_8_9_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_9_10_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_8_10_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_8_10_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_8_10_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_8_10_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_8_10_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_8_10_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_8_10_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_8_10_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_8_10_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_8_10_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_8_10_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_8_10_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_7_10_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_8_11_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_8_9_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_9_10_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_7_10_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_8_11_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_8_9_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_9_10_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_7_10_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_8_11_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_8_9_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_9_10_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_8_10_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_8_10_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_8_10_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_8_10_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_8_10_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_8_10_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_8_10_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_8_10_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_8_10_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_8_10_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_8_10_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_8_10_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_7_10_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_8_11_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_8_9_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_9_10_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_7_10_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_8_11_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_8_9_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_9_10_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_7_10_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_8_11_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_8_9_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_9_10_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_8_10_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_8_10_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_8_10_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_8_10_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_8_10_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_8_10_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_8_10_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_8_10_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_8_10_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_8_10_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_8_10_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_8_10_out_S_noc3_yummy )
);


tile
tile154 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[154] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd10),
    .default_coreid_y           (8'd9),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd154)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[154]   )
    ,.unavailable_o       ( unavailable_o[154] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[154]   )
    ,.ipi_i               ( ipi_i[154]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[154*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile154_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile154_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_8_10_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_9_11_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_9_9_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_10_10_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_8_10_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_9_11_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_9_9_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_10_10_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_8_10_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_9_11_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_9_9_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_10_10_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_9_10_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_9_10_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_9_10_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_9_10_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_9_10_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_9_10_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_9_10_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_9_10_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_9_10_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_9_10_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_9_10_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_9_10_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_8_10_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_9_11_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_9_9_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_10_10_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_8_10_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_9_11_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_9_9_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_10_10_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_8_10_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_9_11_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_9_9_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_10_10_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_9_10_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_9_10_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_9_10_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_9_10_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_9_10_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_9_10_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_9_10_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_9_10_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_9_10_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_9_10_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_9_10_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_9_10_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_8_10_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_9_11_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_9_9_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_10_10_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_8_10_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_9_11_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_9_9_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_10_10_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_8_10_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_9_11_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_9_9_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_10_10_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_9_10_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_9_10_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_9_10_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_9_10_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_9_10_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_9_10_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_9_10_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_9_10_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_9_10_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_9_10_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_9_10_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_9_10_out_S_noc3_yummy )
);


tile
tile170 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[170] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd10),
    .default_coreid_y           (8'd10),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd170)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[170]   )
    ,.unavailable_o       ( unavailable_o[170] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[170]   )
    ,.ipi_i               ( ipi_i[170]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[170*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile170_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile170_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_9_10_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_10_11_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_10_9_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_11_10_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_9_10_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_10_11_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_10_9_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_11_10_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_9_10_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_10_11_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_10_9_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_11_10_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_10_10_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_10_10_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_10_10_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_10_10_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_10_10_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_10_10_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_10_10_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_10_10_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_10_10_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_10_10_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_10_10_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_10_10_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_9_10_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_10_11_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_10_9_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_11_10_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_9_10_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_10_11_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_10_9_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_11_10_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_9_10_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_10_11_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_10_9_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_11_10_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_10_10_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_10_10_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_10_10_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_10_10_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_10_10_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_10_10_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_10_10_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_10_10_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_10_10_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_10_10_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_10_10_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_10_10_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_9_10_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_10_11_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_10_9_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_11_10_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_9_10_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_10_11_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_10_9_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_11_10_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_9_10_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_10_11_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_10_9_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_11_10_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_10_10_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_10_10_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_10_10_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_10_10_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_10_10_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_10_10_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_10_10_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_10_10_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_10_10_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_10_10_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_10_10_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_10_10_out_S_noc3_yummy )
);


tile
tile186 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[186] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd10),
    .default_coreid_y           (8'd11),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd186)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[186]   )
    ,.unavailable_o       ( unavailable_o[186] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[186]   )
    ,.ipi_i               ( ipi_i[186]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[186*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile186_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile186_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_10_10_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_11_11_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_11_9_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_12_10_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_10_10_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_11_11_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_11_9_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_12_10_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_10_10_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_11_11_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_11_9_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_12_10_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_11_10_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_11_10_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_11_10_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_11_10_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_11_10_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_11_10_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_11_10_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_11_10_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_11_10_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_11_10_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_11_10_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_11_10_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_10_10_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_11_11_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_11_9_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_12_10_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_10_10_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_11_11_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_11_9_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_12_10_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_10_10_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_11_11_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_11_9_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_12_10_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_11_10_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_11_10_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_11_10_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_11_10_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_11_10_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_11_10_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_11_10_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_11_10_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_11_10_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_11_10_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_11_10_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_11_10_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_10_10_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_11_11_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_11_9_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_12_10_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_10_10_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_11_11_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_11_9_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_12_10_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_10_10_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_11_11_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_11_9_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_12_10_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_11_10_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_11_10_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_11_10_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_11_10_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_11_10_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_11_10_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_11_10_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_11_10_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_11_10_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_11_10_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_11_10_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_11_10_out_S_noc3_yummy )
);


tile
tile202 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[202] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd10),
    .default_coreid_y           (8'd12),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd202)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[202]   )
    ,.unavailable_o       ( unavailable_o[202] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[202]   )
    ,.ipi_i               ( ipi_i[202]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[202*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile202_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile202_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_11_10_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_12_11_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_12_9_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_13_10_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_11_10_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_12_11_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_12_9_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_13_10_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_11_10_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_12_11_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_12_9_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_13_10_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_12_10_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_12_10_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_12_10_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_12_10_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_12_10_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_12_10_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_12_10_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_12_10_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_12_10_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_12_10_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_12_10_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_12_10_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_11_10_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_12_11_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_12_9_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_13_10_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_11_10_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_12_11_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_12_9_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_13_10_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_11_10_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_12_11_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_12_9_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_13_10_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_12_10_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_12_10_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_12_10_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_12_10_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_12_10_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_12_10_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_12_10_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_12_10_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_12_10_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_12_10_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_12_10_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_12_10_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_11_10_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_12_11_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_12_9_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_13_10_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_11_10_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_12_11_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_12_9_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_13_10_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_11_10_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_12_11_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_12_9_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_13_10_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_12_10_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_12_10_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_12_10_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_12_10_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_12_10_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_12_10_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_12_10_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_12_10_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_12_10_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_12_10_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_12_10_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_12_10_out_S_noc3_yummy )
);


tile
tile218 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[218] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd10),
    .default_coreid_y           (8'd13),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd218)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[218]   )
    ,.unavailable_o       ( unavailable_o[218] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[218]   )
    ,.ipi_i               ( ipi_i[218]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[218*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile218_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile218_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_12_10_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_13_11_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_13_9_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_14_10_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_12_10_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_13_11_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_13_9_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_14_10_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_12_10_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_13_11_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_13_9_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_14_10_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_13_10_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_13_10_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_13_10_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_13_10_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_13_10_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_13_10_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_13_10_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_13_10_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_13_10_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_13_10_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_13_10_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_13_10_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_12_10_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_13_11_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_13_9_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_14_10_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_12_10_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_13_11_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_13_9_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_14_10_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_12_10_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_13_11_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_13_9_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_14_10_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_13_10_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_13_10_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_13_10_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_13_10_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_13_10_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_13_10_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_13_10_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_13_10_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_13_10_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_13_10_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_13_10_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_13_10_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_12_10_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_13_11_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_13_9_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_14_10_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_12_10_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_13_11_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_13_9_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_14_10_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_12_10_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_13_11_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_13_9_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_14_10_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_13_10_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_13_10_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_13_10_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_13_10_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_13_10_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_13_10_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_13_10_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_13_10_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_13_10_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_13_10_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_13_10_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_13_10_out_S_noc3_yummy )
);


tile
tile234 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[234] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd10),
    .default_coreid_y           (8'd14),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd234)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[234]   )
    ,.unavailable_o       ( unavailable_o[234] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[234]   )
    ,.ipi_i               ( ipi_i[234]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[234*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile234_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile234_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_13_10_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_14_11_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_14_9_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_15_10_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_13_10_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_14_11_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_14_9_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_15_10_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_13_10_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_14_11_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_14_9_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_15_10_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_14_10_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_14_10_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_14_10_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_14_10_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_14_10_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_14_10_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_14_10_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_14_10_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_14_10_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_14_10_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_14_10_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_14_10_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_13_10_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_14_11_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_14_9_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_15_10_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_13_10_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_14_11_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_14_9_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_15_10_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_13_10_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_14_11_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_14_9_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_15_10_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_14_10_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_14_10_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_14_10_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_14_10_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_14_10_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_14_10_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_14_10_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_14_10_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_14_10_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_14_10_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_14_10_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_14_10_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_13_10_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_14_11_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_14_9_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_15_10_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_13_10_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_14_11_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_14_9_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_15_10_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_13_10_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_14_11_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_14_9_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_15_10_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_14_10_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_14_10_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_14_10_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_14_10_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_14_10_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_14_10_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_14_10_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_14_10_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_14_10_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_14_10_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_14_10_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_14_10_out_S_noc3_yummy )
);


tile
tile250 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[250] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd10),
    .default_coreid_y           (8'd15),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd250)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[250]   )
    ,.unavailable_o       ( unavailable_o[250] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[250]   )
    ,.ipi_i               ( ipi_i[250]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[250*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile250_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile250_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_14_10_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_15_11_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_15_9_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( dummy_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_14_10_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_15_11_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_15_9_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( dummy_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_14_10_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_15_11_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_15_9_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( dummy_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_15_10_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_15_10_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_15_10_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_15_10_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_15_10_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_15_10_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_15_10_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_15_10_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_15_10_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_15_10_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_15_10_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_15_10_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_14_10_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_15_11_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_15_9_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( dummy_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_14_10_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_15_11_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_15_9_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( dummy_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_14_10_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_15_11_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_15_9_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( dummy_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_15_10_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_15_10_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_15_10_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_15_10_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_15_10_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_15_10_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_15_10_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_15_10_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_15_10_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_15_10_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_15_10_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_15_10_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_14_10_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_15_11_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_15_9_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( dummy_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_14_10_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_15_11_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_15_9_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( dummy_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_14_10_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_15_11_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_15_9_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( dummy_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_15_10_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_15_10_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_15_10_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_15_10_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_15_10_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_15_10_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_15_10_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_15_10_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_15_10_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_15_10_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_15_10_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_15_10_out_S_noc3_yummy )
);


tile
tile11 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[11] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd11),
    .default_coreid_y           (8'd0),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd11)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[11]   )
    ,.unavailable_o       ( unavailable_o[11] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[11]   )
    ,.ipi_i               ( ipi_i[11]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[11*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile11_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile11_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( dummy_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_0_12_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_0_10_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_1_11_out_N_noc1_data   ),
    .dyn0_validIn_N      ( dummy_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_0_12_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_0_10_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_1_11_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( dummy_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_0_12_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_0_10_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_1_11_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_0_11_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_0_11_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_0_11_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_0_11_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_0_11_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_0_11_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_0_11_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_0_11_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_0_11_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_0_11_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_0_11_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_0_11_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( dummy_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_0_12_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_0_10_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_1_11_out_N_noc2_data   ),
    .dyn1_validIn_N      ( dummy_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_0_12_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_0_10_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_1_11_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( dummy_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_0_12_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_0_10_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_1_11_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_0_11_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_0_11_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_0_11_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_0_11_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_0_11_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_0_11_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_0_11_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_0_11_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_0_11_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_0_11_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_0_11_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_0_11_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( dummy_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_0_12_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_0_10_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_1_11_out_N_noc3_data   ),
    .dyn2_validIn_N      ( dummy_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_0_12_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_0_10_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_1_11_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( dummy_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_0_12_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_0_10_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_1_11_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_0_11_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_0_11_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_0_11_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_0_11_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_0_11_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_0_11_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_0_11_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_0_11_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_0_11_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_0_11_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_0_11_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_0_11_out_S_noc3_yummy )
);


tile
tile27 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[27] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd11),
    .default_coreid_y           (8'd1),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd27)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[27]   )
    ,.unavailable_o       ( unavailable_o[27] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[27]   )
    ,.ipi_i               ( ipi_i[27]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[27*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile27_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile27_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_0_11_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_1_12_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_1_10_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_2_11_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_0_11_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_1_12_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_1_10_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_2_11_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_0_11_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_1_12_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_1_10_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_2_11_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_1_11_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_1_11_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_1_11_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_1_11_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_1_11_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_1_11_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_1_11_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_1_11_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_1_11_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_1_11_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_1_11_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_1_11_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_0_11_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_1_12_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_1_10_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_2_11_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_0_11_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_1_12_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_1_10_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_2_11_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_0_11_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_1_12_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_1_10_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_2_11_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_1_11_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_1_11_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_1_11_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_1_11_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_1_11_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_1_11_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_1_11_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_1_11_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_1_11_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_1_11_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_1_11_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_1_11_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_0_11_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_1_12_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_1_10_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_2_11_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_0_11_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_1_12_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_1_10_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_2_11_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_0_11_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_1_12_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_1_10_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_2_11_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_1_11_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_1_11_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_1_11_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_1_11_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_1_11_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_1_11_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_1_11_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_1_11_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_1_11_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_1_11_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_1_11_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_1_11_out_S_noc3_yummy )
);


tile
tile43 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[43] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd11),
    .default_coreid_y           (8'd2),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd43)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[43]   )
    ,.unavailable_o       ( unavailable_o[43] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[43]   )
    ,.ipi_i               ( ipi_i[43]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[43*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile43_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile43_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_1_11_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_2_12_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_2_10_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_3_11_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_1_11_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_2_12_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_2_10_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_3_11_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_1_11_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_2_12_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_2_10_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_3_11_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_2_11_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_2_11_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_2_11_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_2_11_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_2_11_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_2_11_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_2_11_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_2_11_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_2_11_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_2_11_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_2_11_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_2_11_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_1_11_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_2_12_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_2_10_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_3_11_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_1_11_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_2_12_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_2_10_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_3_11_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_1_11_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_2_12_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_2_10_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_3_11_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_2_11_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_2_11_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_2_11_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_2_11_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_2_11_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_2_11_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_2_11_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_2_11_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_2_11_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_2_11_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_2_11_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_2_11_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_1_11_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_2_12_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_2_10_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_3_11_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_1_11_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_2_12_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_2_10_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_3_11_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_1_11_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_2_12_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_2_10_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_3_11_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_2_11_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_2_11_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_2_11_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_2_11_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_2_11_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_2_11_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_2_11_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_2_11_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_2_11_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_2_11_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_2_11_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_2_11_out_S_noc3_yummy )
);


tile
tile59 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[59] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd11),
    .default_coreid_y           (8'd3),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd59)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[59]   )
    ,.unavailable_o       ( unavailable_o[59] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[59]   )
    ,.ipi_i               ( ipi_i[59]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[59*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile59_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile59_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_2_11_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_3_12_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_3_10_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_4_11_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_2_11_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_3_12_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_3_10_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_4_11_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_2_11_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_3_12_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_3_10_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_4_11_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_3_11_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_3_11_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_3_11_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_3_11_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_3_11_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_3_11_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_3_11_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_3_11_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_3_11_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_3_11_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_3_11_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_3_11_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_2_11_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_3_12_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_3_10_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_4_11_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_2_11_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_3_12_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_3_10_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_4_11_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_2_11_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_3_12_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_3_10_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_4_11_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_3_11_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_3_11_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_3_11_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_3_11_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_3_11_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_3_11_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_3_11_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_3_11_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_3_11_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_3_11_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_3_11_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_3_11_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_2_11_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_3_12_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_3_10_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_4_11_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_2_11_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_3_12_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_3_10_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_4_11_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_2_11_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_3_12_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_3_10_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_4_11_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_3_11_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_3_11_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_3_11_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_3_11_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_3_11_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_3_11_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_3_11_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_3_11_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_3_11_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_3_11_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_3_11_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_3_11_out_S_noc3_yummy )
);


tile
tile75 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[75] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd11),
    .default_coreid_y           (8'd4),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd75)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[75]   )
    ,.unavailable_o       ( unavailable_o[75] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[75]   )
    ,.ipi_i               ( ipi_i[75]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[75*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile75_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile75_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_3_11_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_4_12_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_4_10_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_5_11_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_3_11_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_4_12_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_4_10_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_5_11_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_3_11_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_4_12_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_4_10_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_5_11_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_4_11_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_4_11_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_4_11_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_4_11_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_4_11_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_4_11_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_4_11_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_4_11_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_4_11_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_4_11_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_4_11_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_4_11_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_3_11_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_4_12_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_4_10_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_5_11_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_3_11_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_4_12_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_4_10_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_5_11_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_3_11_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_4_12_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_4_10_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_5_11_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_4_11_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_4_11_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_4_11_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_4_11_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_4_11_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_4_11_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_4_11_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_4_11_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_4_11_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_4_11_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_4_11_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_4_11_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_3_11_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_4_12_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_4_10_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_5_11_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_3_11_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_4_12_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_4_10_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_5_11_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_3_11_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_4_12_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_4_10_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_5_11_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_4_11_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_4_11_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_4_11_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_4_11_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_4_11_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_4_11_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_4_11_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_4_11_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_4_11_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_4_11_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_4_11_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_4_11_out_S_noc3_yummy )
);


tile
tile91 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[91] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd11),
    .default_coreid_y           (8'd5),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd91)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[91]   )
    ,.unavailable_o       ( unavailable_o[91] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[91]   )
    ,.ipi_i               ( ipi_i[91]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[91*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile91_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile91_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_4_11_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_5_12_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_5_10_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_6_11_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_4_11_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_5_12_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_5_10_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_6_11_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_4_11_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_5_12_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_5_10_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_6_11_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_5_11_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_5_11_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_5_11_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_5_11_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_5_11_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_5_11_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_5_11_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_5_11_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_5_11_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_5_11_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_5_11_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_5_11_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_4_11_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_5_12_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_5_10_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_6_11_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_4_11_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_5_12_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_5_10_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_6_11_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_4_11_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_5_12_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_5_10_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_6_11_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_5_11_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_5_11_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_5_11_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_5_11_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_5_11_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_5_11_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_5_11_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_5_11_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_5_11_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_5_11_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_5_11_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_5_11_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_4_11_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_5_12_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_5_10_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_6_11_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_4_11_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_5_12_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_5_10_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_6_11_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_4_11_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_5_12_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_5_10_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_6_11_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_5_11_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_5_11_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_5_11_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_5_11_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_5_11_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_5_11_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_5_11_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_5_11_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_5_11_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_5_11_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_5_11_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_5_11_out_S_noc3_yummy )
);


tile
tile107 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[107] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd11),
    .default_coreid_y           (8'd6),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd107)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[107]   )
    ,.unavailable_o       ( unavailable_o[107] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[107]   )
    ,.ipi_i               ( ipi_i[107]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[107*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile107_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile107_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_5_11_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_6_12_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_6_10_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_7_11_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_5_11_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_6_12_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_6_10_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_7_11_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_5_11_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_6_12_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_6_10_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_7_11_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_6_11_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_6_11_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_6_11_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_6_11_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_6_11_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_6_11_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_6_11_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_6_11_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_6_11_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_6_11_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_6_11_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_6_11_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_5_11_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_6_12_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_6_10_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_7_11_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_5_11_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_6_12_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_6_10_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_7_11_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_5_11_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_6_12_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_6_10_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_7_11_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_6_11_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_6_11_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_6_11_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_6_11_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_6_11_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_6_11_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_6_11_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_6_11_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_6_11_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_6_11_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_6_11_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_6_11_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_5_11_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_6_12_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_6_10_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_7_11_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_5_11_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_6_12_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_6_10_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_7_11_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_5_11_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_6_12_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_6_10_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_7_11_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_6_11_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_6_11_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_6_11_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_6_11_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_6_11_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_6_11_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_6_11_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_6_11_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_6_11_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_6_11_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_6_11_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_6_11_out_S_noc3_yummy )
);


tile
tile123 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[123] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd11),
    .default_coreid_y           (8'd7),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd123)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[123]   )
    ,.unavailable_o       ( unavailable_o[123] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[123]   )
    ,.ipi_i               ( ipi_i[123]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[123*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile123_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile123_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_6_11_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_7_12_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_7_10_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_8_11_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_6_11_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_7_12_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_7_10_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_8_11_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_6_11_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_7_12_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_7_10_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_8_11_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_7_11_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_7_11_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_7_11_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_7_11_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_7_11_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_7_11_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_7_11_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_7_11_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_7_11_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_7_11_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_7_11_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_7_11_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_6_11_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_7_12_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_7_10_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_8_11_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_6_11_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_7_12_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_7_10_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_8_11_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_6_11_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_7_12_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_7_10_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_8_11_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_7_11_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_7_11_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_7_11_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_7_11_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_7_11_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_7_11_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_7_11_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_7_11_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_7_11_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_7_11_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_7_11_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_7_11_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_6_11_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_7_12_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_7_10_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_8_11_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_6_11_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_7_12_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_7_10_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_8_11_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_6_11_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_7_12_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_7_10_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_8_11_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_7_11_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_7_11_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_7_11_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_7_11_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_7_11_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_7_11_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_7_11_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_7_11_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_7_11_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_7_11_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_7_11_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_7_11_out_S_noc3_yummy )
);


tile
tile139 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[139] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd11),
    .default_coreid_y           (8'd8),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd139)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[139]   )
    ,.unavailable_o       ( unavailable_o[139] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[139]   )
    ,.ipi_i               ( ipi_i[139]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[139*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile139_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile139_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_7_11_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_8_12_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_8_10_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_9_11_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_7_11_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_8_12_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_8_10_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_9_11_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_7_11_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_8_12_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_8_10_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_9_11_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_8_11_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_8_11_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_8_11_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_8_11_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_8_11_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_8_11_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_8_11_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_8_11_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_8_11_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_8_11_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_8_11_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_8_11_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_7_11_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_8_12_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_8_10_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_9_11_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_7_11_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_8_12_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_8_10_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_9_11_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_7_11_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_8_12_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_8_10_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_9_11_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_8_11_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_8_11_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_8_11_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_8_11_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_8_11_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_8_11_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_8_11_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_8_11_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_8_11_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_8_11_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_8_11_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_8_11_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_7_11_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_8_12_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_8_10_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_9_11_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_7_11_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_8_12_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_8_10_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_9_11_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_7_11_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_8_12_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_8_10_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_9_11_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_8_11_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_8_11_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_8_11_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_8_11_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_8_11_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_8_11_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_8_11_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_8_11_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_8_11_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_8_11_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_8_11_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_8_11_out_S_noc3_yummy )
);


tile
tile155 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[155] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd11),
    .default_coreid_y           (8'd9),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd155)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[155]   )
    ,.unavailable_o       ( unavailable_o[155] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[155]   )
    ,.ipi_i               ( ipi_i[155]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[155*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile155_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile155_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_8_11_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_9_12_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_9_10_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_10_11_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_8_11_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_9_12_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_9_10_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_10_11_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_8_11_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_9_12_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_9_10_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_10_11_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_9_11_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_9_11_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_9_11_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_9_11_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_9_11_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_9_11_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_9_11_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_9_11_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_9_11_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_9_11_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_9_11_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_9_11_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_8_11_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_9_12_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_9_10_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_10_11_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_8_11_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_9_12_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_9_10_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_10_11_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_8_11_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_9_12_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_9_10_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_10_11_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_9_11_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_9_11_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_9_11_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_9_11_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_9_11_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_9_11_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_9_11_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_9_11_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_9_11_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_9_11_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_9_11_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_9_11_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_8_11_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_9_12_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_9_10_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_10_11_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_8_11_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_9_12_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_9_10_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_10_11_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_8_11_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_9_12_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_9_10_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_10_11_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_9_11_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_9_11_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_9_11_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_9_11_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_9_11_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_9_11_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_9_11_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_9_11_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_9_11_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_9_11_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_9_11_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_9_11_out_S_noc3_yummy )
);


tile
tile171 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[171] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd11),
    .default_coreid_y           (8'd10),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd171)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[171]   )
    ,.unavailable_o       ( unavailable_o[171] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[171]   )
    ,.ipi_i               ( ipi_i[171]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[171*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile171_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile171_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_9_11_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_10_12_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_10_10_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_11_11_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_9_11_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_10_12_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_10_10_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_11_11_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_9_11_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_10_12_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_10_10_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_11_11_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_10_11_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_10_11_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_10_11_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_10_11_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_10_11_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_10_11_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_10_11_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_10_11_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_10_11_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_10_11_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_10_11_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_10_11_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_9_11_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_10_12_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_10_10_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_11_11_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_9_11_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_10_12_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_10_10_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_11_11_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_9_11_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_10_12_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_10_10_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_11_11_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_10_11_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_10_11_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_10_11_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_10_11_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_10_11_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_10_11_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_10_11_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_10_11_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_10_11_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_10_11_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_10_11_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_10_11_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_9_11_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_10_12_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_10_10_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_11_11_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_9_11_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_10_12_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_10_10_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_11_11_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_9_11_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_10_12_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_10_10_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_11_11_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_10_11_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_10_11_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_10_11_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_10_11_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_10_11_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_10_11_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_10_11_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_10_11_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_10_11_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_10_11_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_10_11_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_10_11_out_S_noc3_yummy )
);


tile
tile187 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[187] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd11),
    .default_coreid_y           (8'd11),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd187)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[187]   )
    ,.unavailable_o       ( unavailable_o[187] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[187]   )
    ,.ipi_i               ( ipi_i[187]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[187*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile187_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile187_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_10_11_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_11_12_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_11_10_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_12_11_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_10_11_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_11_12_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_11_10_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_12_11_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_10_11_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_11_12_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_11_10_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_12_11_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_11_11_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_11_11_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_11_11_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_11_11_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_11_11_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_11_11_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_11_11_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_11_11_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_11_11_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_11_11_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_11_11_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_11_11_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_10_11_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_11_12_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_11_10_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_12_11_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_10_11_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_11_12_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_11_10_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_12_11_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_10_11_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_11_12_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_11_10_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_12_11_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_11_11_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_11_11_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_11_11_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_11_11_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_11_11_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_11_11_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_11_11_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_11_11_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_11_11_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_11_11_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_11_11_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_11_11_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_10_11_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_11_12_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_11_10_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_12_11_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_10_11_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_11_12_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_11_10_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_12_11_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_10_11_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_11_12_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_11_10_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_12_11_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_11_11_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_11_11_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_11_11_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_11_11_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_11_11_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_11_11_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_11_11_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_11_11_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_11_11_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_11_11_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_11_11_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_11_11_out_S_noc3_yummy )
);


tile
tile203 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[203] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd11),
    .default_coreid_y           (8'd12),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd203)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[203]   )
    ,.unavailable_o       ( unavailable_o[203] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[203]   )
    ,.ipi_i               ( ipi_i[203]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[203*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile203_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile203_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_11_11_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_12_12_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_12_10_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_13_11_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_11_11_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_12_12_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_12_10_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_13_11_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_11_11_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_12_12_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_12_10_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_13_11_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_12_11_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_12_11_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_12_11_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_12_11_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_12_11_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_12_11_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_12_11_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_12_11_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_12_11_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_12_11_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_12_11_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_12_11_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_11_11_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_12_12_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_12_10_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_13_11_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_11_11_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_12_12_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_12_10_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_13_11_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_11_11_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_12_12_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_12_10_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_13_11_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_12_11_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_12_11_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_12_11_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_12_11_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_12_11_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_12_11_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_12_11_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_12_11_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_12_11_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_12_11_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_12_11_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_12_11_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_11_11_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_12_12_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_12_10_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_13_11_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_11_11_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_12_12_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_12_10_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_13_11_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_11_11_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_12_12_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_12_10_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_13_11_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_12_11_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_12_11_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_12_11_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_12_11_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_12_11_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_12_11_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_12_11_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_12_11_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_12_11_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_12_11_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_12_11_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_12_11_out_S_noc3_yummy )
);


tile
tile219 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[219] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd11),
    .default_coreid_y           (8'd13),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd219)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[219]   )
    ,.unavailable_o       ( unavailable_o[219] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[219]   )
    ,.ipi_i               ( ipi_i[219]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[219*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile219_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile219_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_12_11_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_13_12_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_13_10_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_14_11_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_12_11_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_13_12_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_13_10_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_14_11_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_12_11_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_13_12_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_13_10_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_14_11_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_13_11_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_13_11_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_13_11_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_13_11_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_13_11_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_13_11_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_13_11_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_13_11_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_13_11_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_13_11_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_13_11_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_13_11_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_12_11_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_13_12_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_13_10_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_14_11_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_12_11_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_13_12_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_13_10_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_14_11_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_12_11_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_13_12_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_13_10_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_14_11_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_13_11_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_13_11_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_13_11_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_13_11_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_13_11_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_13_11_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_13_11_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_13_11_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_13_11_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_13_11_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_13_11_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_13_11_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_12_11_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_13_12_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_13_10_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_14_11_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_12_11_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_13_12_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_13_10_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_14_11_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_12_11_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_13_12_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_13_10_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_14_11_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_13_11_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_13_11_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_13_11_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_13_11_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_13_11_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_13_11_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_13_11_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_13_11_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_13_11_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_13_11_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_13_11_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_13_11_out_S_noc3_yummy )
);


tile
tile235 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[235] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd11),
    .default_coreid_y           (8'd14),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd235)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[235]   )
    ,.unavailable_o       ( unavailable_o[235] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[235]   )
    ,.ipi_i               ( ipi_i[235]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[235*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile235_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile235_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_13_11_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_14_12_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_14_10_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_15_11_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_13_11_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_14_12_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_14_10_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_15_11_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_13_11_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_14_12_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_14_10_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_15_11_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_14_11_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_14_11_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_14_11_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_14_11_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_14_11_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_14_11_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_14_11_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_14_11_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_14_11_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_14_11_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_14_11_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_14_11_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_13_11_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_14_12_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_14_10_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_15_11_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_13_11_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_14_12_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_14_10_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_15_11_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_13_11_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_14_12_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_14_10_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_15_11_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_14_11_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_14_11_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_14_11_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_14_11_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_14_11_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_14_11_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_14_11_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_14_11_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_14_11_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_14_11_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_14_11_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_14_11_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_13_11_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_14_12_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_14_10_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_15_11_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_13_11_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_14_12_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_14_10_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_15_11_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_13_11_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_14_12_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_14_10_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_15_11_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_14_11_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_14_11_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_14_11_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_14_11_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_14_11_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_14_11_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_14_11_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_14_11_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_14_11_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_14_11_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_14_11_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_14_11_out_S_noc3_yummy )
);


tile
tile251 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[251] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd11),
    .default_coreid_y           (8'd15),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd251)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[251]   )
    ,.unavailable_o       ( unavailable_o[251] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[251]   )
    ,.ipi_i               ( ipi_i[251]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[251*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile251_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile251_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_14_11_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_15_12_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_15_10_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( dummy_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_14_11_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_15_12_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_15_10_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( dummy_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_14_11_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_15_12_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_15_10_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( dummy_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_15_11_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_15_11_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_15_11_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_15_11_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_15_11_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_15_11_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_15_11_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_15_11_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_15_11_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_15_11_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_15_11_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_15_11_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_14_11_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_15_12_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_15_10_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( dummy_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_14_11_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_15_12_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_15_10_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( dummy_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_14_11_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_15_12_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_15_10_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( dummy_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_15_11_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_15_11_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_15_11_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_15_11_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_15_11_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_15_11_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_15_11_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_15_11_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_15_11_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_15_11_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_15_11_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_15_11_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_14_11_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_15_12_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_15_10_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( dummy_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_14_11_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_15_12_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_15_10_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( dummy_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_14_11_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_15_12_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_15_10_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( dummy_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_15_11_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_15_11_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_15_11_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_15_11_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_15_11_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_15_11_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_15_11_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_15_11_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_15_11_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_15_11_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_15_11_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_15_11_out_S_noc3_yummy )
);


tile
tile12 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[12] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd12),
    .default_coreid_y           (8'd0),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd12)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[12]   )
    ,.unavailable_o       ( unavailable_o[12] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[12]   )
    ,.ipi_i               ( ipi_i[12]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[12*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile12_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile12_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( dummy_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_0_13_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_0_11_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_1_12_out_N_noc1_data   ),
    .dyn0_validIn_N      ( dummy_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_0_13_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_0_11_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_1_12_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( dummy_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_0_13_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_0_11_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_1_12_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_0_12_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_0_12_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_0_12_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_0_12_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_0_12_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_0_12_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_0_12_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_0_12_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_0_12_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_0_12_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_0_12_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_0_12_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( dummy_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_0_13_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_0_11_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_1_12_out_N_noc2_data   ),
    .dyn1_validIn_N      ( dummy_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_0_13_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_0_11_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_1_12_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( dummy_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_0_13_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_0_11_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_1_12_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_0_12_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_0_12_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_0_12_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_0_12_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_0_12_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_0_12_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_0_12_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_0_12_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_0_12_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_0_12_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_0_12_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_0_12_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( dummy_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_0_13_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_0_11_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_1_12_out_N_noc3_data   ),
    .dyn2_validIn_N      ( dummy_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_0_13_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_0_11_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_1_12_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( dummy_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_0_13_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_0_11_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_1_12_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_0_12_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_0_12_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_0_12_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_0_12_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_0_12_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_0_12_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_0_12_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_0_12_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_0_12_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_0_12_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_0_12_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_0_12_out_S_noc3_yummy )
);


tile
tile28 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[28] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd12),
    .default_coreid_y           (8'd1),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd28)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[28]   )
    ,.unavailable_o       ( unavailable_o[28] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[28]   )
    ,.ipi_i               ( ipi_i[28]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[28*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile28_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile28_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_0_12_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_1_13_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_1_11_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_2_12_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_0_12_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_1_13_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_1_11_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_2_12_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_0_12_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_1_13_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_1_11_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_2_12_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_1_12_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_1_12_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_1_12_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_1_12_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_1_12_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_1_12_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_1_12_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_1_12_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_1_12_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_1_12_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_1_12_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_1_12_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_0_12_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_1_13_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_1_11_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_2_12_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_0_12_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_1_13_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_1_11_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_2_12_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_0_12_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_1_13_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_1_11_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_2_12_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_1_12_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_1_12_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_1_12_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_1_12_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_1_12_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_1_12_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_1_12_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_1_12_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_1_12_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_1_12_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_1_12_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_1_12_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_0_12_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_1_13_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_1_11_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_2_12_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_0_12_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_1_13_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_1_11_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_2_12_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_0_12_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_1_13_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_1_11_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_2_12_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_1_12_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_1_12_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_1_12_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_1_12_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_1_12_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_1_12_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_1_12_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_1_12_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_1_12_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_1_12_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_1_12_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_1_12_out_S_noc3_yummy )
);


tile
tile44 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[44] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd12),
    .default_coreid_y           (8'd2),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd44)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[44]   )
    ,.unavailable_o       ( unavailable_o[44] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[44]   )
    ,.ipi_i               ( ipi_i[44]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[44*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile44_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile44_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_1_12_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_2_13_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_2_11_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_3_12_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_1_12_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_2_13_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_2_11_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_3_12_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_1_12_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_2_13_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_2_11_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_3_12_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_2_12_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_2_12_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_2_12_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_2_12_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_2_12_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_2_12_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_2_12_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_2_12_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_2_12_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_2_12_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_2_12_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_2_12_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_1_12_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_2_13_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_2_11_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_3_12_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_1_12_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_2_13_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_2_11_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_3_12_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_1_12_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_2_13_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_2_11_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_3_12_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_2_12_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_2_12_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_2_12_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_2_12_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_2_12_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_2_12_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_2_12_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_2_12_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_2_12_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_2_12_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_2_12_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_2_12_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_1_12_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_2_13_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_2_11_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_3_12_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_1_12_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_2_13_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_2_11_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_3_12_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_1_12_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_2_13_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_2_11_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_3_12_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_2_12_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_2_12_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_2_12_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_2_12_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_2_12_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_2_12_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_2_12_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_2_12_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_2_12_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_2_12_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_2_12_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_2_12_out_S_noc3_yummy )
);


tile
tile60 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[60] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd12),
    .default_coreid_y           (8'd3),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd60)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[60]   )
    ,.unavailable_o       ( unavailable_o[60] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[60]   )
    ,.ipi_i               ( ipi_i[60]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[60*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile60_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile60_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_2_12_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_3_13_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_3_11_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_4_12_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_2_12_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_3_13_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_3_11_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_4_12_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_2_12_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_3_13_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_3_11_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_4_12_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_3_12_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_3_12_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_3_12_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_3_12_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_3_12_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_3_12_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_3_12_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_3_12_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_3_12_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_3_12_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_3_12_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_3_12_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_2_12_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_3_13_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_3_11_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_4_12_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_2_12_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_3_13_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_3_11_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_4_12_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_2_12_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_3_13_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_3_11_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_4_12_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_3_12_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_3_12_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_3_12_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_3_12_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_3_12_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_3_12_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_3_12_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_3_12_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_3_12_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_3_12_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_3_12_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_3_12_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_2_12_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_3_13_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_3_11_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_4_12_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_2_12_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_3_13_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_3_11_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_4_12_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_2_12_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_3_13_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_3_11_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_4_12_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_3_12_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_3_12_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_3_12_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_3_12_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_3_12_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_3_12_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_3_12_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_3_12_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_3_12_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_3_12_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_3_12_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_3_12_out_S_noc3_yummy )
);


tile
tile76 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[76] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd12),
    .default_coreid_y           (8'd4),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd76)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[76]   )
    ,.unavailable_o       ( unavailable_o[76] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[76]   )
    ,.ipi_i               ( ipi_i[76]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[76*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile76_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile76_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_3_12_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_4_13_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_4_11_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_5_12_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_3_12_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_4_13_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_4_11_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_5_12_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_3_12_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_4_13_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_4_11_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_5_12_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_4_12_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_4_12_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_4_12_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_4_12_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_4_12_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_4_12_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_4_12_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_4_12_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_4_12_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_4_12_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_4_12_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_4_12_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_3_12_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_4_13_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_4_11_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_5_12_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_3_12_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_4_13_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_4_11_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_5_12_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_3_12_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_4_13_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_4_11_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_5_12_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_4_12_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_4_12_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_4_12_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_4_12_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_4_12_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_4_12_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_4_12_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_4_12_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_4_12_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_4_12_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_4_12_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_4_12_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_3_12_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_4_13_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_4_11_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_5_12_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_3_12_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_4_13_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_4_11_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_5_12_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_3_12_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_4_13_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_4_11_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_5_12_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_4_12_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_4_12_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_4_12_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_4_12_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_4_12_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_4_12_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_4_12_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_4_12_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_4_12_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_4_12_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_4_12_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_4_12_out_S_noc3_yummy )
);


tile
tile92 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[92] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd12),
    .default_coreid_y           (8'd5),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd92)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[92]   )
    ,.unavailable_o       ( unavailable_o[92] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[92]   )
    ,.ipi_i               ( ipi_i[92]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[92*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile92_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile92_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_4_12_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_5_13_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_5_11_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_6_12_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_4_12_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_5_13_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_5_11_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_6_12_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_4_12_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_5_13_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_5_11_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_6_12_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_5_12_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_5_12_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_5_12_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_5_12_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_5_12_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_5_12_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_5_12_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_5_12_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_5_12_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_5_12_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_5_12_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_5_12_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_4_12_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_5_13_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_5_11_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_6_12_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_4_12_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_5_13_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_5_11_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_6_12_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_4_12_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_5_13_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_5_11_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_6_12_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_5_12_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_5_12_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_5_12_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_5_12_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_5_12_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_5_12_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_5_12_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_5_12_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_5_12_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_5_12_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_5_12_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_5_12_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_4_12_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_5_13_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_5_11_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_6_12_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_4_12_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_5_13_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_5_11_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_6_12_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_4_12_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_5_13_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_5_11_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_6_12_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_5_12_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_5_12_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_5_12_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_5_12_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_5_12_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_5_12_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_5_12_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_5_12_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_5_12_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_5_12_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_5_12_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_5_12_out_S_noc3_yummy )
);


tile
tile108 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[108] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd12),
    .default_coreid_y           (8'd6),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd108)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[108]   )
    ,.unavailable_o       ( unavailable_o[108] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[108]   )
    ,.ipi_i               ( ipi_i[108]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[108*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile108_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile108_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_5_12_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_6_13_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_6_11_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_7_12_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_5_12_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_6_13_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_6_11_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_7_12_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_5_12_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_6_13_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_6_11_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_7_12_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_6_12_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_6_12_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_6_12_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_6_12_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_6_12_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_6_12_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_6_12_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_6_12_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_6_12_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_6_12_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_6_12_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_6_12_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_5_12_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_6_13_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_6_11_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_7_12_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_5_12_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_6_13_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_6_11_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_7_12_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_5_12_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_6_13_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_6_11_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_7_12_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_6_12_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_6_12_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_6_12_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_6_12_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_6_12_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_6_12_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_6_12_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_6_12_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_6_12_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_6_12_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_6_12_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_6_12_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_5_12_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_6_13_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_6_11_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_7_12_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_5_12_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_6_13_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_6_11_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_7_12_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_5_12_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_6_13_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_6_11_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_7_12_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_6_12_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_6_12_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_6_12_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_6_12_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_6_12_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_6_12_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_6_12_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_6_12_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_6_12_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_6_12_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_6_12_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_6_12_out_S_noc3_yummy )
);


tile
tile124 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[124] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd12),
    .default_coreid_y           (8'd7),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd124)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[124]   )
    ,.unavailable_o       ( unavailable_o[124] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[124]   )
    ,.ipi_i               ( ipi_i[124]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[124*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile124_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile124_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_6_12_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_7_13_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_7_11_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_8_12_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_6_12_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_7_13_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_7_11_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_8_12_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_6_12_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_7_13_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_7_11_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_8_12_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_7_12_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_7_12_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_7_12_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_7_12_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_7_12_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_7_12_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_7_12_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_7_12_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_7_12_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_7_12_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_7_12_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_7_12_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_6_12_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_7_13_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_7_11_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_8_12_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_6_12_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_7_13_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_7_11_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_8_12_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_6_12_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_7_13_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_7_11_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_8_12_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_7_12_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_7_12_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_7_12_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_7_12_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_7_12_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_7_12_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_7_12_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_7_12_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_7_12_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_7_12_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_7_12_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_7_12_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_6_12_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_7_13_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_7_11_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_8_12_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_6_12_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_7_13_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_7_11_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_8_12_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_6_12_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_7_13_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_7_11_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_8_12_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_7_12_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_7_12_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_7_12_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_7_12_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_7_12_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_7_12_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_7_12_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_7_12_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_7_12_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_7_12_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_7_12_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_7_12_out_S_noc3_yummy )
);


tile
tile140 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[140] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd12),
    .default_coreid_y           (8'd8),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd140)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[140]   )
    ,.unavailable_o       ( unavailable_o[140] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[140]   )
    ,.ipi_i               ( ipi_i[140]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[140*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile140_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile140_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_7_12_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_8_13_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_8_11_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_9_12_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_7_12_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_8_13_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_8_11_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_9_12_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_7_12_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_8_13_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_8_11_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_9_12_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_8_12_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_8_12_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_8_12_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_8_12_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_8_12_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_8_12_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_8_12_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_8_12_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_8_12_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_8_12_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_8_12_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_8_12_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_7_12_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_8_13_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_8_11_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_9_12_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_7_12_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_8_13_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_8_11_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_9_12_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_7_12_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_8_13_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_8_11_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_9_12_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_8_12_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_8_12_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_8_12_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_8_12_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_8_12_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_8_12_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_8_12_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_8_12_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_8_12_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_8_12_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_8_12_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_8_12_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_7_12_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_8_13_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_8_11_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_9_12_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_7_12_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_8_13_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_8_11_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_9_12_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_7_12_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_8_13_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_8_11_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_9_12_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_8_12_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_8_12_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_8_12_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_8_12_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_8_12_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_8_12_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_8_12_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_8_12_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_8_12_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_8_12_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_8_12_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_8_12_out_S_noc3_yummy )
);


tile
tile156 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[156] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd12),
    .default_coreid_y           (8'd9),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd156)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[156]   )
    ,.unavailable_o       ( unavailable_o[156] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[156]   )
    ,.ipi_i               ( ipi_i[156]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[156*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile156_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile156_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_8_12_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_9_13_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_9_11_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_10_12_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_8_12_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_9_13_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_9_11_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_10_12_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_8_12_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_9_13_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_9_11_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_10_12_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_9_12_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_9_12_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_9_12_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_9_12_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_9_12_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_9_12_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_9_12_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_9_12_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_9_12_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_9_12_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_9_12_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_9_12_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_8_12_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_9_13_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_9_11_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_10_12_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_8_12_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_9_13_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_9_11_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_10_12_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_8_12_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_9_13_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_9_11_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_10_12_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_9_12_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_9_12_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_9_12_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_9_12_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_9_12_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_9_12_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_9_12_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_9_12_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_9_12_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_9_12_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_9_12_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_9_12_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_8_12_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_9_13_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_9_11_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_10_12_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_8_12_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_9_13_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_9_11_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_10_12_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_8_12_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_9_13_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_9_11_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_10_12_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_9_12_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_9_12_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_9_12_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_9_12_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_9_12_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_9_12_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_9_12_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_9_12_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_9_12_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_9_12_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_9_12_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_9_12_out_S_noc3_yummy )
);


tile
tile172 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[172] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd12),
    .default_coreid_y           (8'd10),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd172)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[172]   )
    ,.unavailable_o       ( unavailable_o[172] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[172]   )
    ,.ipi_i               ( ipi_i[172]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[172*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile172_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile172_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_9_12_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_10_13_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_10_11_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_11_12_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_9_12_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_10_13_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_10_11_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_11_12_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_9_12_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_10_13_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_10_11_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_11_12_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_10_12_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_10_12_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_10_12_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_10_12_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_10_12_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_10_12_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_10_12_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_10_12_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_10_12_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_10_12_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_10_12_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_10_12_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_9_12_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_10_13_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_10_11_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_11_12_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_9_12_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_10_13_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_10_11_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_11_12_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_9_12_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_10_13_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_10_11_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_11_12_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_10_12_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_10_12_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_10_12_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_10_12_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_10_12_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_10_12_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_10_12_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_10_12_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_10_12_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_10_12_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_10_12_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_10_12_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_9_12_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_10_13_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_10_11_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_11_12_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_9_12_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_10_13_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_10_11_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_11_12_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_9_12_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_10_13_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_10_11_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_11_12_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_10_12_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_10_12_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_10_12_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_10_12_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_10_12_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_10_12_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_10_12_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_10_12_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_10_12_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_10_12_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_10_12_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_10_12_out_S_noc3_yummy )
);


tile
tile188 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[188] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd12),
    .default_coreid_y           (8'd11),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd188)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[188]   )
    ,.unavailable_o       ( unavailable_o[188] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[188]   )
    ,.ipi_i               ( ipi_i[188]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[188*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile188_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile188_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_10_12_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_11_13_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_11_11_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_12_12_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_10_12_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_11_13_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_11_11_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_12_12_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_10_12_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_11_13_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_11_11_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_12_12_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_11_12_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_11_12_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_11_12_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_11_12_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_11_12_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_11_12_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_11_12_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_11_12_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_11_12_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_11_12_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_11_12_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_11_12_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_10_12_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_11_13_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_11_11_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_12_12_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_10_12_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_11_13_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_11_11_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_12_12_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_10_12_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_11_13_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_11_11_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_12_12_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_11_12_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_11_12_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_11_12_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_11_12_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_11_12_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_11_12_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_11_12_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_11_12_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_11_12_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_11_12_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_11_12_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_11_12_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_10_12_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_11_13_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_11_11_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_12_12_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_10_12_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_11_13_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_11_11_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_12_12_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_10_12_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_11_13_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_11_11_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_12_12_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_11_12_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_11_12_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_11_12_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_11_12_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_11_12_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_11_12_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_11_12_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_11_12_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_11_12_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_11_12_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_11_12_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_11_12_out_S_noc3_yummy )
);


tile
tile204 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[204] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd12),
    .default_coreid_y           (8'd12),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd204)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[204]   )
    ,.unavailable_o       ( unavailable_o[204] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[204]   )
    ,.ipi_i               ( ipi_i[204]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[204*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile204_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile204_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_11_12_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_12_13_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_12_11_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_13_12_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_11_12_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_12_13_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_12_11_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_13_12_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_11_12_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_12_13_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_12_11_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_13_12_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_12_12_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_12_12_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_12_12_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_12_12_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_12_12_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_12_12_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_12_12_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_12_12_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_12_12_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_12_12_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_12_12_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_12_12_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_11_12_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_12_13_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_12_11_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_13_12_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_11_12_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_12_13_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_12_11_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_13_12_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_11_12_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_12_13_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_12_11_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_13_12_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_12_12_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_12_12_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_12_12_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_12_12_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_12_12_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_12_12_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_12_12_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_12_12_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_12_12_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_12_12_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_12_12_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_12_12_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_11_12_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_12_13_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_12_11_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_13_12_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_11_12_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_12_13_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_12_11_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_13_12_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_11_12_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_12_13_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_12_11_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_13_12_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_12_12_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_12_12_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_12_12_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_12_12_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_12_12_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_12_12_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_12_12_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_12_12_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_12_12_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_12_12_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_12_12_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_12_12_out_S_noc3_yummy )
);


tile
tile220 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[220] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd12),
    .default_coreid_y           (8'd13),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd220)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[220]   )
    ,.unavailable_o       ( unavailable_o[220] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[220]   )
    ,.ipi_i               ( ipi_i[220]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[220*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile220_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile220_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_12_12_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_13_13_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_13_11_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_14_12_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_12_12_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_13_13_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_13_11_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_14_12_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_12_12_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_13_13_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_13_11_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_14_12_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_13_12_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_13_12_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_13_12_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_13_12_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_13_12_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_13_12_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_13_12_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_13_12_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_13_12_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_13_12_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_13_12_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_13_12_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_12_12_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_13_13_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_13_11_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_14_12_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_12_12_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_13_13_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_13_11_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_14_12_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_12_12_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_13_13_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_13_11_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_14_12_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_13_12_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_13_12_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_13_12_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_13_12_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_13_12_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_13_12_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_13_12_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_13_12_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_13_12_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_13_12_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_13_12_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_13_12_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_12_12_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_13_13_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_13_11_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_14_12_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_12_12_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_13_13_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_13_11_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_14_12_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_12_12_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_13_13_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_13_11_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_14_12_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_13_12_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_13_12_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_13_12_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_13_12_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_13_12_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_13_12_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_13_12_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_13_12_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_13_12_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_13_12_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_13_12_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_13_12_out_S_noc3_yummy )
);


tile
tile236 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[236] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd12),
    .default_coreid_y           (8'd14),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd236)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[236]   )
    ,.unavailable_o       ( unavailable_o[236] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[236]   )
    ,.ipi_i               ( ipi_i[236]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[236*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile236_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile236_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_13_12_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_14_13_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_14_11_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_15_12_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_13_12_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_14_13_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_14_11_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_15_12_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_13_12_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_14_13_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_14_11_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_15_12_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_14_12_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_14_12_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_14_12_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_14_12_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_14_12_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_14_12_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_14_12_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_14_12_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_14_12_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_14_12_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_14_12_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_14_12_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_13_12_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_14_13_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_14_11_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_15_12_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_13_12_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_14_13_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_14_11_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_15_12_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_13_12_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_14_13_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_14_11_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_15_12_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_14_12_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_14_12_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_14_12_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_14_12_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_14_12_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_14_12_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_14_12_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_14_12_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_14_12_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_14_12_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_14_12_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_14_12_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_13_12_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_14_13_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_14_11_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_15_12_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_13_12_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_14_13_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_14_11_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_15_12_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_13_12_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_14_13_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_14_11_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_15_12_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_14_12_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_14_12_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_14_12_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_14_12_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_14_12_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_14_12_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_14_12_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_14_12_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_14_12_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_14_12_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_14_12_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_14_12_out_S_noc3_yummy )
);


tile
tile252 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[252] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd12),
    .default_coreid_y           (8'd15),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd252)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[252]   )
    ,.unavailable_o       ( unavailable_o[252] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[252]   )
    ,.ipi_i               ( ipi_i[252]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[252*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile252_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile252_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_14_12_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_15_13_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_15_11_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( dummy_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_14_12_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_15_13_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_15_11_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( dummy_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_14_12_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_15_13_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_15_11_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( dummy_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_15_12_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_15_12_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_15_12_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_15_12_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_15_12_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_15_12_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_15_12_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_15_12_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_15_12_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_15_12_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_15_12_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_15_12_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_14_12_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_15_13_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_15_11_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( dummy_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_14_12_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_15_13_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_15_11_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( dummy_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_14_12_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_15_13_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_15_11_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( dummy_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_15_12_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_15_12_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_15_12_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_15_12_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_15_12_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_15_12_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_15_12_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_15_12_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_15_12_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_15_12_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_15_12_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_15_12_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_14_12_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_15_13_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_15_11_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( dummy_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_14_12_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_15_13_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_15_11_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( dummy_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_14_12_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_15_13_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_15_11_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( dummy_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_15_12_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_15_12_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_15_12_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_15_12_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_15_12_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_15_12_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_15_12_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_15_12_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_15_12_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_15_12_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_15_12_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_15_12_out_S_noc3_yummy )
);


tile
tile13 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[13] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd13),
    .default_coreid_y           (8'd0),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd13)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[13]   )
    ,.unavailable_o       ( unavailable_o[13] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[13]   )
    ,.ipi_i               ( ipi_i[13]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[13*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile13_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile13_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( dummy_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_0_14_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_0_12_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_1_13_out_N_noc1_data   ),
    .dyn0_validIn_N      ( dummy_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_0_14_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_0_12_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_1_13_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( dummy_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_0_14_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_0_12_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_1_13_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_0_13_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_0_13_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_0_13_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_0_13_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_0_13_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_0_13_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_0_13_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_0_13_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_0_13_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_0_13_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_0_13_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_0_13_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( dummy_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_0_14_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_0_12_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_1_13_out_N_noc2_data   ),
    .dyn1_validIn_N      ( dummy_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_0_14_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_0_12_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_1_13_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( dummy_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_0_14_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_0_12_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_1_13_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_0_13_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_0_13_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_0_13_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_0_13_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_0_13_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_0_13_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_0_13_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_0_13_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_0_13_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_0_13_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_0_13_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_0_13_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( dummy_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_0_14_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_0_12_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_1_13_out_N_noc3_data   ),
    .dyn2_validIn_N      ( dummy_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_0_14_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_0_12_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_1_13_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( dummy_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_0_14_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_0_12_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_1_13_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_0_13_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_0_13_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_0_13_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_0_13_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_0_13_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_0_13_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_0_13_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_0_13_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_0_13_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_0_13_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_0_13_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_0_13_out_S_noc3_yummy )
);


tile
tile29 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[29] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd13),
    .default_coreid_y           (8'd1),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd29)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[29]   )
    ,.unavailable_o       ( unavailable_o[29] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[29]   )
    ,.ipi_i               ( ipi_i[29]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[29*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile29_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile29_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_0_13_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_1_14_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_1_12_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_2_13_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_0_13_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_1_14_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_1_12_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_2_13_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_0_13_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_1_14_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_1_12_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_2_13_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_1_13_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_1_13_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_1_13_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_1_13_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_1_13_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_1_13_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_1_13_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_1_13_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_1_13_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_1_13_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_1_13_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_1_13_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_0_13_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_1_14_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_1_12_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_2_13_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_0_13_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_1_14_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_1_12_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_2_13_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_0_13_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_1_14_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_1_12_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_2_13_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_1_13_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_1_13_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_1_13_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_1_13_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_1_13_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_1_13_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_1_13_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_1_13_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_1_13_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_1_13_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_1_13_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_1_13_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_0_13_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_1_14_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_1_12_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_2_13_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_0_13_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_1_14_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_1_12_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_2_13_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_0_13_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_1_14_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_1_12_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_2_13_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_1_13_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_1_13_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_1_13_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_1_13_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_1_13_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_1_13_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_1_13_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_1_13_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_1_13_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_1_13_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_1_13_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_1_13_out_S_noc3_yummy )
);


tile
tile45 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[45] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd13),
    .default_coreid_y           (8'd2),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd45)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[45]   )
    ,.unavailable_o       ( unavailable_o[45] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[45]   )
    ,.ipi_i               ( ipi_i[45]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[45*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile45_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile45_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_1_13_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_2_14_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_2_12_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_3_13_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_1_13_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_2_14_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_2_12_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_3_13_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_1_13_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_2_14_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_2_12_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_3_13_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_2_13_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_2_13_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_2_13_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_2_13_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_2_13_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_2_13_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_2_13_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_2_13_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_2_13_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_2_13_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_2_13_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_2_13_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_1_13_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_2_14_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_2_12_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_3_13_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_1_13_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_2_14_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_2_12_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_3_13_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_1_13_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_2_14_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_2_12_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_3_13_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_2_13_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_2_13_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_2_13_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_2_13_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_2_13_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_2_13_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_2_13_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_2_13_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_2_13_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_2_13_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_2_13_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_2_13_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_1_13_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_2_14_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_2_12_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_3_13_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_1_13_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_2_14_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_2_12_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_3_13_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_1_13_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_2_14_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_2_12_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_3_13_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_2_13_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_2_13_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_2_13_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_2_13_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_2_13_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_2_13_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_2_13_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_2_13_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_2_13_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_2_13_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_2_13_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_2_13_out_S_noc3_yummy )
);


tile
tile61 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[61] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd13),
    .default_coreid_y           (8'd3),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd61)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[61]   )
    ,.unavailable_o       ( unavailable_o[61] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[61]   )
    ,.ipi_i               ( ipi_i[61]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[61*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile61_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile61_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_2_13_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_3_14_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_3_12_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_4_13_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_2_13_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_3_14_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_3_12_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_4_13_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_2_13_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_3_14_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_3_12_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_4_13_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_3_13_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_3_13_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_3_13_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_3_13_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_3_13_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_3_13_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_3_13_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_3_13_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_3_13_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_3_13_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_3_13_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_3_13_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_2_13_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_3_14_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_3_12_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_4_13_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_2_13_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_3_14_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_3_12_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_4_13_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_2_13_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_3_14_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_3_12_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_4_13_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_3_13_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_3_13_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_3_13_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_3_13_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_3_13_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_3_13_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_3_13_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_3_13_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_3_13_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_3_13_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_3_13_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_3_13_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_2_13_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_3_14_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_3_12_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_4_13_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_2_13_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_3_14_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_3_12_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_4_13_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_2_13_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_3_14_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_3_12_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_4_13_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_3_13_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_3_13_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_3_13_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_3_13_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_3_13_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_3_13_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_3_13_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_3_13_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_3_13_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_3_13_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_3_13_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_3_13_out_S_noc3_yummy )
);


tile
tile77 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[77] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd13),
    .default_coreid_y           (8'd4),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd77)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[77]   )
    ,.unavailable_o       ( unavailable_o[77] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[77]   )
    ,.ipi_i               ( ipi_i[77]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[77*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile77_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile77_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_3_13_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_4_14_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_4_12_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_5_13_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_3_13_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_4_14_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_4_12_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_5_13_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_3_13_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_4_14_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_4_12_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_5_13_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_4_13_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_4_13_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_4_13_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_4_13_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_4_13_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_4_13_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_4_13_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_4_13_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_4_13_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_4_13_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_4_13_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_4_13_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_3_13_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_4_14_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_4_12_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_5_13_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_3_13_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_4_14_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_4_12_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_5_13_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_3_13_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_4_14_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_4_12_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_5_13_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_4_13_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_4_13_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_4_13_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_4_13_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_4_13_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_4_13_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_4_13_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_4_13_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_4_13_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_4_13_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_4_13_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_4_13_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_3_13_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_4_14_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_4_12_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_5_13_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_3_13_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_4_14_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_4_12_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_5_13_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_3_13_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_4_14_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_4_12_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_5_13_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_4_13_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_4_13_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_4_13_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_4_13_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_4_13_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_4_13_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_4_13_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_4_13_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_4_13_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_4_13_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_4_13_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_4_13_out_S_noc3_yummy )
);


tile
tile93 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[93] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd13),
    .default_coreid_y           (8'd5),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd93)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[93]   )
    ,.unavailable_o       ( unavailable_o[93] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[93]   )
    ,.ipi_i               ( ipi_i[93]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[93*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile93_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile93_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_4_13_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_5_14_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_5_12_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_6_13_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_4_13_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_5_14_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_5_12_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_6_13_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_4_13_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_5_14_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_5_12_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_6_13_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_5_13_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_5_13_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_5_13_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_5_13_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_5_13_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_5_13_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_5_13_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_5_13_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_5_13_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_5_13_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_5_13_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_5_13_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_4_13_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_5_14_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_5_12_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_6_13_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_4_13_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_5_14_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_5_12_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_6_13_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_4_13_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_5_14_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_5_12_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_6_13_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_5_13_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_5_13_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_5_13_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_5_13_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_5_13_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_5_13_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_5_13_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_5_13_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_5_13_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_5_13_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_5_13_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_5_13_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_4_13_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_5_14_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_5_12_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_6_13_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_4_13_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_5_14_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_5_12_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_6_13_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_4_13_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_5_14_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_5_12_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_6_13_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_5_13_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_5_13_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_5_13_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_5_13_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_5_13_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_5_13_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_5_13_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_5_13_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_5_13_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_5_13_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_5_13_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_5_13_out_S_noc3_yummy )
);


tile
tile109 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[109] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd13),
    .default_coreid_y           (8'd6),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd109)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[109]   )
    ,.unavailable_o       ( unavailable_o[109] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[109]   )
    ,.ipi_i               ( ipi_i[109]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[109*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile109_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile109_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_5_13_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_6_14_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_6_12_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_7_13_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_5_13_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_6_14_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_6_12_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_7_13_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_5_13_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_6_14_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_6_12_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_7_13_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_6_13_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_6_13_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_6_13_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_6_13_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_6_13_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_6_13_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_6_13_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_6_13_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_6_13_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_6_13_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_6_13_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_6_13_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_5_13_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_6_14_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_6_12_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_7_13_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_5_13_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_6_14_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_6_12_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_7_13_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_5_13_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_6_14_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_6_12_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_7_13_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_6_13_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_6_13_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_6_13_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_6_13_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_6_13_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_6_13_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_6_13_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_6_13_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_6_13_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_6_13_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_6_13_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_6_13_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_5_13_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_6_14_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_6_12_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_7_13_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_5_13_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_6_14_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_6_12_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_7_13_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_5_13_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_6_14_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_6_12_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_7_13_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_6_13_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_6_13_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_6_13_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_6_13_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_6_13_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_6_13_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_6_13_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_6_13_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_6_13_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_6_13_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_6_13_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_6_13_out_S_noc3_yummy )
);


tile
tile125 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[125] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd13),
    .default_coreid_y           (8'd7),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd125)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[125]   )
    ,.unavailable_o       ( unavailable_o[125] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[125]   )
    ,.ipi_i               ( ipi_i[125]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[125*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile125_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile125_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_6_13_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_7_14_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_7_12_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_8_13_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_6_13_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_7_14_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_7_12_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_8_13_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_6_13_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_7_14_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_7_12_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_8_13_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_7_13_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_7_13_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_7_13_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_7_13_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_7_13_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_7_13_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_7_13_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_7_13_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_7_13_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_7_13_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_7_13_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_7_13_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_6_13_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_7_14_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_7_12_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_8_13_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_6_13_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_7_14_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_7_12_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_8_13_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_6_13_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_7_14_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_7_12_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_8_13_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_7_13_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_7_13_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_7_13_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_7_13_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_7_13_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_7_13_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_7_13_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_7_13_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_7_13_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_7_13_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_7_13_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_7_13_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_6_13_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_7_14_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_7_12_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_8_13_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_6_13_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_7_14_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_7_12_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_8_13_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_6_13_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_7_14_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_7_12_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_8_13_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_7_13_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_7_13_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_7_13_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_7_13_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_7_13_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_7_13_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_7_13_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_7_13_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_7_13_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_7_13_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_7_13_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_7_13_out_S_noc3_yummy )
);


tile
tile141 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[141] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd13),
    .default_coreid_y           (8'd8),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd141)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[141]   )
    ,.unavailable_o       ( unavailable_o[141] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[141]   )
    ,.ipi_i               ( ipi_i[141]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[141*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile141_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile141_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_7_13_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_8_14_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_8_12_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_9_13_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_7_13_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_8_14_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_8_12_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_9_13_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_7_13_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_8_14_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_8_12_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_9_13_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_8_13_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_8_13_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_8_13_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_8_13_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_8_13_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_8_13_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_8_13_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_8_13_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_8_13_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_8_13_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_8_13_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_8_13_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_7_13_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_8_14_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_8_12_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_9_13_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_7_13_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_8_14_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_8_12_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_9_13_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_7_13_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_8_14_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_8_12_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_9_13_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_8_13_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_8_13_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_8_13_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_8_13_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_8_13_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_8_13_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_8_13_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_8_13_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_8_13_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_8_13_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_8_13_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_8_13_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_7_13_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_8_14_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_8_12_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_9_13_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_7_13_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_8_14_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_8_12_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_9_13_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_7_13_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_8_14_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_8_12_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_9_13_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_8_13_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_8_13_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_8_13_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_8_13_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_8_13_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_8_13_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_8_13_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_8_13_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_8_13_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_8_13_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_8_13_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_8_13_out_S_noc3_yummy )
);


tile
tile157 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[157] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd13),
    .default_coreid_y           (8'd9),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd157)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[157]   )
    ,.unavailable_o       ( unavailable_o[157] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[157]   )
    ,.ipi_i               ( ipi_i[157]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[157*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile157_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile157_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_8_13_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_9_14_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_9_12_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_10_13_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_8_13_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_9_14_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_9_12_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_10_13_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_8_13_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_9_14_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_9_12_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_10_13_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_9_13_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_9_13_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_9_13_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_9_13_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_9_13_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_9_13_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_9_13_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_9_13_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_9_13_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_9_13_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_9_13_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_9_13_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_8_13_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_9_14_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_9_12_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_10_13_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_8_13_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_9_14_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_9_12_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_10_13_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_8_13_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_9_14_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_9_12_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_10_13_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_9_13_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_9_13_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_9_13_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_9_13_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_9_13_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_9_13_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_9_13_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_9_13_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_9_13_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_9_13_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_9_13_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_9_13_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_8_13_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_9_14_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_9_12_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_10_13_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_8_13_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_9_14_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_9_12_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_10_13_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_8_13_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_9_14_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_9_12_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_10_13_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_9_13_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_9_13_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_9_13_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_9_13_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_9_13_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_9_13_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_9_13_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_9_13_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_9_13_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_9_13_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_9_13_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_9_13_out_S_noc3_yummy )
);


tile
tile173 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[173] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd13),
    .default_coreid_y           (8'd10),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd173)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[173]   )
    ,.unavailable_o       ( unavailable_o[173] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[173]   )
    ,.ipi_i               ( ipi_i[173]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[173*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile173_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile173_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_9_13_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_10_14_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_10_12_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_11_13_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_9_13_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_10_14_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_10_12_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_11_13_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_9_13_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_10_14_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_10_12_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_11_13_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_10_13_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_10_13_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_10_13_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_10_13_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_10_13_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_10_13_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_10_13_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_10_13_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_10_13_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_10_13_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_10_13_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_10_13_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_9_13_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_10_14_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_10_12_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_11_13_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_9_13_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_10_14_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_10_12_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_11_13_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_9_13_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_10_14_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_10_12_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_11_13_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_10_13_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_10_13_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_10_13_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_10_13_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_10_13_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_10_13_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_10_13_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_10_13_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_10_13_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_10_13_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_10_13_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_10_13_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_9_13_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_10_14_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_10_12_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_11_13_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_9_13_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_10_14_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_10_12_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_11_13_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_9_13_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_10_14_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_10_12_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_11_13_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_10_13_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_10_13_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_10_13_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_10_13_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_10_13_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_10_13_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_10_13_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_10_13_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_10_13_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_10_13_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_10_13_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_10_13_out_S_noc3_yummy )
);


tile
tile189 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[189] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd13),
    .default_coreid_y           (8'd11),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd189)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[189]   )
    ,.unavailable_o       ( unavailable_o[189] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[189]   )
    ,.ipi_i               ( ipi_i[189]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[189*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile189_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile189_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_10_13_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_11_14_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_11_12_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_12_13_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_10_13_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_11_14_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_11_12_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_12_13_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_10_13_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_11_14_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_11_12_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_12_13_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_11_13_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_11_13_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_11_13_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_11_13_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_11_13_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_11_13_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_11_13_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_11_13_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_11_13_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_11_13_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_11_13_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_11_13_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_10_13_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_11_14_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_11_12_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_12_13_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_10_13_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_11_14_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_11_12_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_12_13_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_10_13_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_11_14_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_11_12_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_12_13_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_11_13_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_11_13_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_11_13_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_11_13_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_11_13_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_11_13_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_11_13_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_11_13_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_11_13_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_11_13_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_11_13_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_11_13_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_10_13_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_11_14_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_11_12_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_12_13_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_10_13_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_11_14_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_11_12_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_12_13_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_10_13_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_11_14_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_11_12_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_12_13_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_11_13_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_11_13_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_11_13_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_11_13_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_11_13_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_11_13_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_11_13_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_11_13_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_11_13_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_11_13_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_11_13_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_11_13_out_S_noc3_yummy )
);


tile
tile205 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[205] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd13),
    .default_coreid_y           (8'd12),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd205)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[205]   )
    ,.unavailable_o       ( unavailable_o[205] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[205]   )
    ,.ipi_i               ( ipi_i[205]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[205*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile205_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile205_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_11_13_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_12_14_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_12_12_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_13_13_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_11_13_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_12_14_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_12_12_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_13_13_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_11_13_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_12_14_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_12_12_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_13_13_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_12_13_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_12_13_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_12_13_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_12_13_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_12_13_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_12_13_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_12_13_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_12_13_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_12_13_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_12_13_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_12_13_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_12_13_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_11_13_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_12_14_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_12_12_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_13_13_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_11_13_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_12_14_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_12_12_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_13_13_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_11_13_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_12_14_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_12_12_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_13_13_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_12_13_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_12_13_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_12_13_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_12_13_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_12_13_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_12_13_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_12_13_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_12_13_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_12_13_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_12_13_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_12_13_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_12_13_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_11_13_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_12_14_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_12_12_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_13_13_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_11_13_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_12_14_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_12_12_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_13_13_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_11_13_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_12_14_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_12_12_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_13_13_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_12_13_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_12_13_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_12_13_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_12_13_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_12_13_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_12_13_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_12_13_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_12_13_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_12_13_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_12_13_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_12_13_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_12_13_out_S_noc3_yummy )
);


tile
tile221 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[221] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd13),
    .default_coreid_y           (8'd13),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd221)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[221]   )
    ,.unavailable_o       ( unavailable_o[221] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[221]   )
    ,.ipi_i               ( ipi_i[221]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[221*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile221_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile221_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_12_13_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_13_14_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_13_12_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_14_13_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_12_13_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_13_14_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_13_12_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_14_13_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_12_13_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_13_14_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_13_12_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_14_13_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_13_13_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_13_13_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_13_13_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_13_13_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_13_13_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_13_13_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_13_13_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_13_13_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_13_13_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_13_13_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_13_13_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_13_13_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_12_13_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_13_14_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_13_12_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_14_13_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_12_13_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_13_14_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_13_12_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_14_13_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_12_13_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_13_14_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_13_12_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_14_13_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_13_13_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_13_13_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_13_13_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_13_13_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_13_13_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_13_13_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_13_13_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_13_13_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_13_13_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_13_13_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_13_13_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_13_13_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_12_13_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_13_14_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_13_12_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_14_13_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_12_13_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_13_14_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_13_12_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_14_13_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_12_13_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_13_14_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_13_12_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_14_13_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_13_13_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_13_13_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_13_13_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_13_13_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_13_13_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_13_13_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_13_13_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_13_13_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_13_13_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_13_13_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_13_13_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_13_13_out_S_noc3_yummy )
);


tile
tile237 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[237] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd13),
    .default_coreid_y           (8'd14),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd237)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[237]   )
    ,.unavailable_o       ( unavailable_o[237] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[237]   )
    ,.ipi_i               ( ipi_i[237]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[237*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile237_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile237_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_13_13_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_14_14_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_14_12_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_15_13_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_13_13_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_14_14_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_14_12_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_15_13_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_13_13_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_14_14_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_14_12_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_15_13_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_14_13_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_14_13_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_14_13_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_14_13_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_14_13_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_14_13_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_14_13_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_14_13_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_14_13_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_14_13_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_14_13_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_14_13_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_13_13_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_14_14_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_14_12_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_15_13_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_13_13_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_14_14_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_14_12_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_15_13_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_13_13_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_14_14_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_14_12_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_15_13_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_14_13_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_14_13_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_14_13_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_14_13_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_14_13_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_14_13_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_14_13_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_14_13_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_14_13_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_14_13_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_14_13_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_14_13_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_13_13_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_14_14_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_14_12_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_15_13_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_13_13_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_14_14_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_14_12_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_15_13_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_13_13_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_14_14_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_14_12_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_15_13_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_14_13_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_14_13_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_14_13_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_14_13_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_14_13_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_14_13_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_14_13_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_14_13_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_14_13_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_14_13_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_14_13_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_14_13_out_S_noc3_yummy )
);


tile
tile253 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[253] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd13),
    .default_coreid_y           (8'd15),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd253)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[253]   )
    ,.unavailable_o       ( unavailable_o[253] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[253]   )
    ,.ipi_i               ( ipi_i[253]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[253*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile253_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile253_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_14_13_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_15_14_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_15_12_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( dummy_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_14_13_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_15_14_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_15_12_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( dummy_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_14_13_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_15_14_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_15_12_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( dummy_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_15_13_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_15_13_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_15_13_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_15_13_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_15_13_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_15_13_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_15_13_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_15_13_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_15_13_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_15_13_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_15_13_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_15_13_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_14_13_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_15_14_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_15_12_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( dummy_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_14_13_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_15_14_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_15_12_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( dummy_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_14_13_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_15_14_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_15_12_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( dummy_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_15_13_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_15_13_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_15_13_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_15_13_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_15_13_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_15_13_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_15_13_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_15_13_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_15_13_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_15_13_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_15_13_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_15_13_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_14_13_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_15_14_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_15_12_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( dummy_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_14_13_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_15_14_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_15_12_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( dummy_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_14_13_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_15_14_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_15_12_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( dummy_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_15_13_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_15_13_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_15_13_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_15_13_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_15_13_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_15_13_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_15_13_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_15_13_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_15_13_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_15_13_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_15_13_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_15_13_out_S_noc3_yummy )
);


tile
tile14 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[14] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd14),
    .default_coreid_y           (8'd0),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd14)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[14]   )
    ,.unavailable_o       ( unavailable_o[14] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[14]   )
    ,.ipi_i               ( ipi_i[14]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[14*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile14_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile14_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( dummy_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_0_15_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_0_13_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_1_14_out_N_noc1_data   ),
    .dyn0_validIn_N      ( dummy_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_0_15_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_0_13_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_1_14_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( dummy_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_0_15_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_0_13_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_1_14_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_0_14_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_0_14_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_0_14_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_0_14_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_0_14_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_0_14_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_0_14_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_0_14_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_0_14_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_0_14_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_0_14_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_0_14_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( dummy_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_0_15_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_0_13_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_1_14_out_N_noc2_data   ),
    .dyn1_validIn_N      ( dummy_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_0_15_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_0_13_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_1_14_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( dummy_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_0_15_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_0_13_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_1_14_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_0_14_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_0_14_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_0_14_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_0_14_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_0_14_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_0_14_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_0_14_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_0_14_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_0_14_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_0_14_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_0_14_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_0_14_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( dummy_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_0_15_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_0_13_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_1_14_out_N_noc3_data   ),
    .dyn2_validIn_N      ( dummy_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_0_15_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_0_13_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_1_14_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( dummy_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_0_15_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_0_13_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_1_14_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_0_14_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_0_14_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_0_14_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_0_14_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_0_14_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_0_14_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_0_14_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_0_14_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_0_14_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_0_14_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_0_14_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_0_14_out_S_noc3_yummy )
);


tile
tile30 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[30] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd14),
    .default_coreid_y           (8'd1),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd30)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[30]   )
    ,.unavailable_o       ( unavailable_o[30] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[30]   )
    ,.ipi_i               ( ipi_i[30]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[30*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile30_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile30_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_0_14_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_1_15_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_1_13_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_2_14_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_0_14_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_1_15_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_1_13_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_2_14_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_0_14_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_1_15_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_1_13_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_2_14_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_1_14_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_1_14_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_1_14_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_1_14_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_1_14_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_1_14_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_1_14_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_1_14_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_1_14_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_1_14_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_1_14_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_1_14_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_0_14_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_1_15_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_1_13_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_2_14_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_0_14_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_1_15_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_1_13_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_2_14_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_0_14_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_1_15_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_1_13_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_2_14_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_1_14_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_1_14_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_1_14_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_1_14_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_1_14_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_1_14_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_1_14_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_1_14_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_1_14_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_1_14_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_1_14_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_1_14_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_0_14_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_1_15_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_1_13_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_2_14_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_0_14_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_1_15_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_1_13_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_2_14_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_0_14_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_1_15_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_1_13_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_2_14_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_1_14_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_1_14_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_1_14_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_1_14_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_1_14_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_1_14_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_1_14_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_1_14_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_1_14_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_1_14_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_1_14_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_1_14_out_S_noc3_yummy )
);


tile
tile46 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[46] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd14),
    .default_coreid_y           (8'd2),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd46)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[46]   )
    ,.unavailable_o       ( unavailable_o[46] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[46]   )
    ,.ipi_i               ( ipi_i[46]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[46*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile46_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile46_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_1_14_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_2_15_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_2_13_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_3_14_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_1_14_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_2_15_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_2_13_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_3_14_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_1_14_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_2_15_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_2_13_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_3_14_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_2_14_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_2_14_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_2_14_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_2_14_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_2_14_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_2_14_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_2_14_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_2_14_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_2_14_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_2_14_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_2_14_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_2_14_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_1_14_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_2_15_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_2_13_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_3_14_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_1_14_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_2_15_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_2_13_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_3_14_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_1_14_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_2_15_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_2_13_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_3_14_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_2_14_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_2_14_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_2_14_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_2_14_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_2_14_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_2_14_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_2_14_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_2_14_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_2_14_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_2_14_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_2_14_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_2_14_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_1_14_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_2_15_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_2_13_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_3_14_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_1_14_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_2_15_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_2_13_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_3_14_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_1_14_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_2_15_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_2_13_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_3_14_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_2_14_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_2_14_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_2_14_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_2_14_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_2_14_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_2_14_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_2_14_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_2_14_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_2_14_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_2_14_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_2_14_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_2_14_out_S_noc3_yummy )
);


tile
tile62 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[62] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd14),
    .default_coreid_y           (8'd3),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd62)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[62]   )
    ,.unavailable_o       ( unavailable_o[62] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[62]   )
    ,.ipi_i               ( ipi_i[62]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[62*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile62_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile62_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_2_14_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_3_15_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_3_13_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_4_14_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_2_14_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_3_15_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_3_13_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_4_14_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_2_14_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_3_15_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_3_13_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_4_14_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_3_14_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_3_14_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_3_14_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_3_14_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_3_14_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_3_14_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_3_14_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_3_14_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_3_14_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_3_14_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_3_14_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_3_14_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_2_14_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_3_15_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_3_13_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_4_14_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_2_14_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_3_15_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_3_13_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_4_14_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_2_14_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_3_15_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_3_13_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_4_14_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_3_14_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_3_14_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_3_14_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_3_14_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_3_14_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_3_14_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_3_14_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_3_14_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_3_14_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_3_14_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_3_14_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_3_14_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_2_14_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_3_15_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_3_13_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_4_14_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_2_14_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_3_15_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_3_13_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_4_14_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_2_14_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_3_15_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_3_13_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_4_14_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_3_14_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_3_14_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_3_14_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_3_14_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_3_14_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_3_14_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_3_14_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_3_14_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_3_14_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_3_14_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_3_14_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_3_14_out_S_noc3_yummy )
);


tile
tile78 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[78] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd14),
    .default_coreid_y           (8'd4),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd78)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[78]   )
    ,.unavailable_o       ( unavailable_o[78] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[78]   )
    ,.ipi_i               ( ipi_i[78]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[78*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile78_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile78_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_3_14_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_4_15_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_4_13_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_5_14_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_3_14_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_4_15_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_4_13_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_5_14_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_3_14_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_4_15_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_4_13_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_5_14_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_4_14_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_4_14_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_4_14_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_4_14_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_4_14_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_4_14_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_4_14_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_4_14_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_4_14_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_4_14_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_4_14_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_4_14_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_3_14_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_4_15_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_4_13_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_5_14_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_3_14_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_4_15_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_4_13_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_5_14_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_3_14_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_4_15_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_4_13_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_5_14_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_4_14_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_4_14_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_4_14_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_4_14_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_4_14_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_4_14_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_4_14_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_4_14_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_4_14_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_4_14_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_4_14_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_4_14_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_3_14_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_4_15_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_4_13_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_5_14_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_3_14_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_4_15_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_4_13_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_5_14_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_3_14_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_4_15_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_4_13_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_5_14_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_4_14_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_4_14_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_4_14_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_4_14_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_4_14_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_4_14_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_4_14_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_4_14_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_4_14_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_4_14_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_4_14_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_4_14_out_S_noc3_yummy )
);


tile
tile94 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[94] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd14),
    .default_coreid_y           (8'd5),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd94)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[94]   )
    ,.unavailable_o       ( unavailable_o[94] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[94]   )
    ,.ipi_i               ( ipi_i[94]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[94*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile94_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile94_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_4_14_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_5_15_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_5_13_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_6_14_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_4_14_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_5_15_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_5_13_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_6_14_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_4_14_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_5_15_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_5_13_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_6_14_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_5_14_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_5_14_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_5_14_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_5_14_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_5_14_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_5_14_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_5_14_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_5_14_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_5_14_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_5_14_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_5_14_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_5_14_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_4_14_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_5_15_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_5_13_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_6_14_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_4_14_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_5_15_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_5_13_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_6_14_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_4_14_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_5_15_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_5_13_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_6_14_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_5_14_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_5_14_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_5_14_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_5_14_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_5_14_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_5_14_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_5_14_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_5_14_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_5_14_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_5_14_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_5_14_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_5_14_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_4_14_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_5_15_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_5_13_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_6_14_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_4_14_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_5_15_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_5_13_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_6_14_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_4_14_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_5_15_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_5_13_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_6_14_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_5_14_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_5_14_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_5_14_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_5_14_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_5_14_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_5_14_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_5_14_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_5_14_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_5_14_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_5_14_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_5_14_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_5_14_out_S_noc3_yummy )
);


tile
tile110 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[110] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd14),
    .default_coreid_y           (8'd6),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd110)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[110]   )
    ,.unavailable_o       ( unavailable_o[110] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[110]   )
    ,.ipi_i               ( ipi_i[110]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[110*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile110_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile110_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_5_14_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_6_15_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_6_13_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_7_14_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_5_14_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_6_15_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_6_13_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_7_14_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_5_14_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_6_15_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_6_13_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_7_14_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_6_14_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_6_14_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_6_14_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_6_14_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_6_14_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_6_14_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_6_14_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_6_14_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_6_14_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_6_14_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_6_14_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_6_14_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_5_14_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_6_15_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_6_13_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_7_14_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_5_14_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_6_15_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_6_13_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_7_14_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_5_14_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_6_15_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_6_13_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_7_14_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_6_14_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_6_14_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_6_14_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_6_14_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_6_14_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_6_14_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_6_14_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_6_14_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_6_14_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_6_14_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_6_14_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_6_14_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_5_14_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_6_15_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_6_13_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_7_14_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_5_14_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_6_15_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_6_13_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_7_14_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_5_14_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_6_15_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_6_13_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_7_14_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_6_14_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_6_14_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_6_14_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_6_14_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_6_14_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_6_14_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_6_14_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_6_14_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_6_14_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_6_14_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_6_14_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_6_14_out_S_noc3_yummy )
);


tile
tile126 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[126] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd14),
    .default_coreid_y           (8'd7),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd126)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[126]   )
    ,.unavailable_o       ( unavailable_o[126] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[126]   )
    ,.ipi_i               ( ipi_i[126]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[126*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile126_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile126_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_6_14_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_7_15_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_7_13_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_8_14_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_6_14_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_7_15_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_7_13_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_8_14_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_6_14_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_7_15_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_7_13_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_8_14_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_7_14_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_7_14_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_7_14_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_7_14_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_7_14_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_7_14_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_7_14_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_7_14_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_7_14_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_7_14_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_7_14_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_7_14_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_6_14_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_7_15_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_7_13_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_8_14_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_6_14_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_7_15_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_7_13_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_8_14_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_6_14_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_7_15_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_7_13_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_8_14_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_7_14_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_7_14_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_7_14_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_7_14_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_7_14_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_7_14_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_7_14_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_7_14_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_7_14_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_7_14_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_7_14_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_7_14_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_6_14_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_7_15_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_7_13_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_8_14_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_6_14_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_7_15_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_7_13_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_8_14_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_6_14_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_7_15_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_7_13_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_8_14_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_7_14_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_7_14_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_7_14_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_7_14_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_7_14_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_7_14_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_7_14_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_7_14_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_7_14_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_7_14_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_7_14_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_7_14_out_S_noc3_yummy )
);


tile
tile142 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[142] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd14),
    .default_coreid_y           (8'd8),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd142)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[142]   )
    ,.unavailable_o       ( unavailable_o[142] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[142]   )
    ,.ipi_i               ( ipi_i[142]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[142*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile142_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile142_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_7_14_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_8_15_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_8_13_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_9_14_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_7_14_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_8_15_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_8_13_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_9_14_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_7_14_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_8_15_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_8_13_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_9_14_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_8_14_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_8_14_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_8_14_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_8_14_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_8_14_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_8_14_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_8_14_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_8_14_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_8_14_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_8_14_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_8_14_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_8_14_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_7_14_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_8_15_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_8_13_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_9_14_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_7_14_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_8_15_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_8_13_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_9_14_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_7_14_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_8_15_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_8_13_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_9_14_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_8_14_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_8_14_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_8_14_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_8_14_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_8_14_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_8_14_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_8_14_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_8_14_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_8_14_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_8_14_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_8_14_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_8_14_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_7_14_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_8_15_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_8_13_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_9_14_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_7_14_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_8_15_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_8_13_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_9_14_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_7_14_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_8_15_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_8_13_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_9_14_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_8_14_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_8_14_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_8_14_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_8_14_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_8_14_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_8_14_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_8_14_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_8_14_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_8_14_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_8_14_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_8_14_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_8_14_out_S_noc3_yummy )
);


tile
tile158 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[158] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd14),
    .default_coreid_y           (8'd9),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd158)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[158]   )
    ,.unavailable_o       ( unavailable_o[158] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[158]   )
    ,.ipi_i               ( ipi_i[158]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[158*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile158_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile158_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_8_14_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_9_15_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_9_13_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_10_14_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_8_14_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_9_15_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_9_13_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_10_14_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_8_14_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_9_15_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_9_13_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_10_14_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_9_14_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_9_14_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_9_14_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_9_14_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_9_14_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_9_14_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_9_14_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_9_14_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_9_14_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_9_14_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_9_14_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_9_14_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_8_14_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_9_15_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_9_13_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_10_14_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_8_14_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_9_15_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_9_13_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_10_14_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_8_14_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_9_15_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_9_13_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_10_14_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_9_14_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_9_14_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_9_14_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_9_14_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_9_14_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_9_14_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_9_14_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_9_14_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_9_14_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_9_14_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_9_14_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_9_14_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_8_14_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_9_15_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_9_13_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_10_14_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_8_14_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_9_15_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_9_13_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_10_14_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_8_14_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_9_15_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_9_13_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_10_14_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_9_14_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_9_14_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_9_14_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_9_14_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_9_14_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_9_14_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_9_14_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_9_14_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_9_14_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_9_14_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_9_14_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_9_14_out_S_noc3_yummy )
);


tile
tile174 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[174] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd14),
    .default_coreid_y           (8'd10),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd174)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[174]   )
    ,.unavailable_o       ( unavailable_o[174] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[174]   )
    ,.ipi_i               ( ipi_i[174]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[174*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile174_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile174_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_9_14_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_10_15_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_10_13_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_11_14_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_9_14_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_10_15_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_10_13_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_11_14_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_9_14_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_10_15_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_10_13_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_11_14_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_10_14_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_10_14_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_10_14_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_10_14_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_10_14_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_10_14_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_10_14_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_10_14_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_10_14_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_10_14_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_10_14_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_10_14_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_9_14_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_10_15_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_10_13_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_11_14_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_9_14_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_10_15_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_10_13_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_11_14_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_9_14_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_10_15_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_10_13_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_11_14_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_10_14_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_10_14_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_10_14_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_10_14_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_10_14_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_10_14_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_10_14_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_10_14_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_10_14_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_10_14_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_10_14_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_10_14_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_9_14_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_10_15_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_10_13_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_11_14_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_9_14_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_10_15_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_10_13_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_11_14_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_9_14_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_10_15_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_10_13_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_11_14_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_10_14_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_10_14_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_10_14_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_10_14_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_10_14_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_10_14_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_10_14_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_10_14_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_10_14_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_10_14_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_10_14_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_10_14_out_S_noc3_yummy )
);


tile
tile190 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[190] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd14),
    .default_coreid_y           (8'd11),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd190)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[190]   )
    ,.unavailable_o       ( unavailable_o[190] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[190]   )
    ,.ipi_i               ( ipi_i[190]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[190*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile190_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile190_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_10_14_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_11_15_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_11_13_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_12_14_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_10_14_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_11_15_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_11_13_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_12_14_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_10_14_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_11_15_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_11_13_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_12_14_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_11_14_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_11_14_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_11_14_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_11_14_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_11_14_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_11_14_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_11_14_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_11_14_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_11_14_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_11_14_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_11_14_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_11_14_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_10_14_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_11_15_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_11_13_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_12_14_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_10_14_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_11_15_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_11_13_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_12_14_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_10_14_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_11_15_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_11_13_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_12_14_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_11_14_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_11_14_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_11_14_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_11_14_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_11_14_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_11_14_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_11_14_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_11_14_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_11_14_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_11_14_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_11_14_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_11_14_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_10_14_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_11_15_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_11_13_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_12_14_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_10_14_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_11_15_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_11_13_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_12_14_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_10_14_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_11_15_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_11_13_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_12_14_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_11_14_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_11_14_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_11_14_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_11_14_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_11_14_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_11_14_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_11_14_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_11_14_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_11_14_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_11_14_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_11_14_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_11_14_out_S_noc3_yummy )
);


tile
tile206 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[206] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd14),
    .default_coreid_y           (8'd12),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd206)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[206]   )
    ,.unavailable_o       ( unavailable_o[206] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[206]   )
    ,.ipi_i               ( ipi_i[206]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[206*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile206_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile206_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_11_14_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_12_15_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_12_13_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_13_14_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_11_14_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_12_15_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_12_13_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_13_14_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_11_14_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_12_15_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_12_13_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_13_14_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_12_14_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_12_14_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_12_14_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_12_14_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_12_14_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_12_14_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_12_14_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_12_14_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_12_14_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_12_14_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_12_14_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_12_14_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_11_14_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_12_15_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_12_13_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_13_14_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_11_14_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_12_15_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_12_13_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_13_14_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_11_14_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_12_15_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_12_13_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_13_14_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_12_14_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_12_14_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_12_14_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_12_14_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_12_14_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_12_14_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_12_14_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_12_14_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_12_14_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_12_14_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_12_14_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_12_14_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_11_14_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_12_15_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_12_13_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_13_14_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_11_14_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_12_15_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_12_13_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_13_14_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_11_14_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_12_15_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_12_13_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_13_14_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_12_14_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_12_14_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_12_14_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_12_14_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_12_14_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_12_14_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_12_14_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_12_14_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_12_14_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_12_14_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_12_14_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_12_14_out_S_noc3_yummy )
);


tile
tile222 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[222] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd14),
    .default_coreid_y           (8'd13),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd222)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[222]   )
    ,.unavailable_o       ( unavailable_o[222] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[222]   )
    ,.ipi_i               ( ipi_i[222]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[222*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile222_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile222_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_12_14_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_13_15_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_13_13_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_14_14_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_12_14_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_13_15_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_13_13_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_14_14_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_12_14_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_13_15_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_13_13_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_14_14_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_13_14_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_13_14_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_13_14_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_13_14_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_13_14_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_13_14_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_13_14_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_13_14_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_13_14_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_13_14_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_13_14_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_13_14_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_12_14_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_13_15_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_13_13_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_14_14_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_12_14_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_13_15_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_13_13_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_14_14_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_12_14_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_13_15_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_13_13_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_14_14_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_13_14_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_13_14_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_13_14_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_13_14_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_13_14_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_13_14_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_13_14_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_13_14_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_13_14_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_13_14_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_13_14_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_13_14_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_12_14_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_13_15_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_13_13_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_14_14_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_12_14_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_13_15_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_13_13_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_14_14_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_12_14_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_13_15_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_13_13_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_14_14_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_13_14_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_13_14_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_13_14_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_13_14_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_13_14_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_13_14_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_13_14_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_13_14_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_13_14_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_13_14_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_13_14_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_13_14_out_S_noc3_yummy )
);


tile
tile238 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[238] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd14),
    .default_coreid_y           (8'd14),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd238)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[238]   )
    ,.unavailable_o       ( unavailable_o[238] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[238]   )
    ,.ipi_i               ( ipi_i[238]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[238*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile238_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile238_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_13_14_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_14_15_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_14_13_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_15_14_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_13_14_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_14_15_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_14_13_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_15_14_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_13_14_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_14_15_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_14_13_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_15_14_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_14_14_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_14_14_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_14_14_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_14_14_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_14_14_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_14_14_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_14_14_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_14_14_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_14_14_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_14_14_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_14_14_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_14_14_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_13_14_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_14_15_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_14_13_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_15_14_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_13_14_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_14_15_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_14_13_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_15_14_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_13_14_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_14_15_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_14_13_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_15_14_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_14_14_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_14_14_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_14_14_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_14_14_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_14_14_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_14_14_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_14_14_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_14_14_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_14_14_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_14_14_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_14_14_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_14_14_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_13_14_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_14_15_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_14_13_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_15_14_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_13_14_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_14_15_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_14_13_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_15_14_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_13_14_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_14_15_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_14_13_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_15_14_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_14_14_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_14_14_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_14_14_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_14_14_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_14_14_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_14_14_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_14_14_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_14_14_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_14_14_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_14_14_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_14_14_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_14_14_out_S_noc3_yummy )
);


tile
tile254 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[254] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd14),
    .default_coreid_y           (8'd15),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd254)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[254]   )
    ,.unavailable_o       ( unavailable_o[254] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[254]   )
    ,.ipi_i               ( ipi_i[254]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[254*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile254_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile254_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_14_14_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( tile_15_15_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_15_13_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( dummy_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_14_14_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( tile_15_15_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_15_13_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( dummy_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_14_14_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( tile_15_15_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_15_13_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( dummy_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_15_14_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_15_14_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_15_14_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_15_14_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_15_14_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_15_14_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_15_14_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_15_14_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_15_14_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_15_14_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_15_14_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_15_14_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_14_14_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( tile_15_15_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_15_13_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( dummy_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_14_14_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( tile_15_15_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_15_13_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( dummy_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_14_14_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( tile_15_15_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_15_13_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( dummy_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_15_14_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_15_14_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_15_14_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_15_14_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_15_14_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_15_14_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_15_14_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_15_14_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_15_14_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_15_14_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_15_14_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_15_14_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_14_14_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( tile_15_15_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_15_13_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( dummy_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_14_14_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( tile_15_15_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_15_13_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( dummy_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_14_14_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( tile_15_15_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_15_13_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( dummy_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_15_14_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_15_14_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_15_14_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_15_14_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_15_14_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_15_14_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_15_14_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_15_14_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_15_14_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_15_14_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_15_14_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_15_14_out_S_noc3_yummy )
);


tile
tile15 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[15] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd15),
    .default_coreid_y           (8'd0),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd15)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[15]   )
    ,.unavailable_o       ( unavailable_o[15] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[15]   )
    ,.ipi_i               ( ipi_i[15]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[15*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile15_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile15_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( dummy_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( dummy_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_0_14_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_1_15_out_N_noc1_data   ),
    .dyn0_validIn_N      ( dummy_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( dummy_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_0_14_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_1_15_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( dummy_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( dummy_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_0_14_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_1_15_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_0_15_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_0_15_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_0_15_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_0_15_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_0_15_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_0_15_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_0_15_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_0_15_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_0_15_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_0_15_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_0_15_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_0_15_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( dummy_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( dummy_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_0_14_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_1_15_out_N_noc2_data   ),
    .dyn1_validIn_N      ( dummy_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( dummy_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_0_14_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_1_15_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( dummy_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( dummy_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_0_14_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_1_15_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_0_15_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_0_15_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_0_15_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_0_15_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_0_15_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_0_15_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_0_15_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_0_15_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_0_15_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_0_15_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_0_15_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_0_15_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( dummy_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( dummy_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_0_14_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_1_15_out_N_noc3_data   ),
    .dyn2_validIn_N      ( dummy_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( dummy_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_0_14_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_1_15_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( dummy_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( dummy_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_0_14_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_1_15_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_0_15_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_0_15_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_0_15_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_0_15_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_0_15_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_0_15_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_0_15_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_0_15_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_0_15_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_0_15_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_0_15_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_0_15_out_S_noc3_yummy )
);


tile
tile31 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[31] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd15),
    .default_coreid_y           (8'd1),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd31)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[31]   )
    ,.unavailable_o       ( unavailable_o[31] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[31]   )
    ,.ipi_i               ( ipi_i[31]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[31*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile31_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile31_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_0_15_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( dummy_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_1_14_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_2_15_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_0_15_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( dummy_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_1_14_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_2_15_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_0_15_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( dummy_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_1_14_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_2_15_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_1_15_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_1_15_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_1_15_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_1_15_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_1_15_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_1_15_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_1_15_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_1_15_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_1_15_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_1_15_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_1_15_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_1_15_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_0_15_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( dummy_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_1_14_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_2_15_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_0_15_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( dummy_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_1_14_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_2_15_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_0_15_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( dummy_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_1_14_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_2_15_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_1_15_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_1_15_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_1_15_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_1_15_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_1_15_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_1_15_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_1_15_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_1_15_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_1_15_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_1_15_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_1_15_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_1_15_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_0_15_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( dummy_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_1_14_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_2_15_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_0_15_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( dummy_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_1_14_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_2_15_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_0_15_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( dummy_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_1_14_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_2_15_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_1_15_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_1_15_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_1_15_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_1_15_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_1_15_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_1_15_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_1_15_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_1_15_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_1_15_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_1_15_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_1_15_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_1_15_out_S_noc3_yummy )
);


tile
tile47 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[47] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd15),
    .default_coreid_y           (8'd2),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd47)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[47]   )
    ,.unavailable_o       ( unavailable_o[47] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[47]   )
    ,.ipi_i               ( ipi_i[47]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[47*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile47_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile47_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_1_15_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( dummy_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_2_14_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_3_15_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_1_15_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( dummy_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_2_14_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_3_15_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_1_15_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( dummy_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_2_14_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_3_15_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_2_15_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_2_15_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_2_15_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_2_15_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_2_15_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_2_15_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_2_15_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_2_15_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_2_15_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_2_15_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_2_15_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_2_15_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_1_15_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( dummy_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_2_14_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_3_15_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_1_15_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( dummy_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_2_14_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_3_15_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_1_15_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( dummy_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_2_14_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_3_15_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_2_15_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_2_15_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_2_15_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_2_15_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_2_15_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_2_15_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_2_15_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_2_15_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_2_15_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_2_15_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_2_15_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_2_15_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_1_15_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( dummy_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_2_14_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_3_15_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_1_15_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( dummy_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_2_14_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_3_15_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_1_15_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( dummy_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_2_14_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_3_15_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_2_15_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_2_15_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_2_15_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_2_15_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_2_15_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_2_15_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_2_15_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_2_15_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_2_15_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_2_15_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_2_15_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_2_15_out_S_noc3_yummy )
);


tile
tile63 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[63] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd15),
    .default_coreid_y           (8'd3),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd63)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[63]   )
    ,.unavailable_o       ( unavailable_o[63] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[63]   )
    ,.ipi_i               ( ipi_i[63]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[63*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile63_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile63_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_2_15_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( dummy_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_3_14_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_4_15_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_2_15_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( dummy_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_3_14_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_4_15_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_2_15_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( dummy_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_3_14_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_4_15_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_3_15_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_3_15_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_3_15_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_3_15_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_3_15_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_3_15_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_3_15_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_3_15_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_3_15_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_3_15_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_3_15_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_3_15_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_2_15_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( dummy_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_3_14_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_4_15_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_2_15_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( dummy_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_3_14_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_4_15_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_2_15_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( dummy_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_3_14_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_4_15_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_3_15_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_3_15_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_3_15_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_3_15_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_3_15_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_3_15_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_3_15_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_3_15_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_3_15_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_3_15_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_3_15_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_3_15_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_2_15_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( dummy_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_3_14_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_4_15_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_2_15_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( dummy_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_3_14_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_4_15_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_2_15_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( dummy_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_3_14_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_4_15_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_3_15_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_3_15_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_3_15_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_3_15_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_3_15_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_3_15_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_3_15_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_3_15_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_3_15_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_3_15_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_3_15_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_3_15_out_S_noc3_yummy )
);


tile
tile79 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[79] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd15),
    .default_coreid_y           (8'd4),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd79)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[79]   )
    ,.unavailable_o       ( unavailable_o[79] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[79]   )
    ,.ipi_i               ( ipi_i[79]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[79*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile79_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile79_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_3_15_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( dummy_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_4_14_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_5_15_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_3_15_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( dummy_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_4_14_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_5_15_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_3_15_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( dummy_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_4_14_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_5_15_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_4_15_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_4_15_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_4_15_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_4_15_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_4_15_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_4_15_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_4_15_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_4_15_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_4_15_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_4_15_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_4_15_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_4_15_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_3_15_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( dummy_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_4_14_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_5_15_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_3_15_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( dummy_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_4_14_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_5_15_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_3_15_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( dummy_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_4_14_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_5_15_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_4_15_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_4_15_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_4_15_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_4_15_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_4_15_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_4_15_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_4_15_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_4_15_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_4_15_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_4_15_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_4_15_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_4_15_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_3_15_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( dummy_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_4_14_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_5_15_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_3_15_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( dummy_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_4_14_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_5_15_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_3_15_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( dummy_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_4_14_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_5_15_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_4_15_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_4_15_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_4_15_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_4_15_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_4_15_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_4_15_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_4_15_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_4_15_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_4_15_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_4_15_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_4_15_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_4_15_out_S_noc3_yummy )
);


tile
tile95 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[95] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd15),
    .default_coreid_y           (8'd5),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd95)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[95]   )
    ,.unavailable_o       ( unavailable_o[95] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[95]   )
    ,.ipi_i               ( ipi_i[95]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[95*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile95_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile95_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_4_15_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( dummy_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_5_14_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_6_15_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_4_15_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( dummy_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_5_14_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_6_15_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_4_15_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( dummy_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_5_14_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_6_15_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_5_15_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_5_15_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_5_15_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_5_15_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_5_15_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_5_15_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_5_15_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_5_15_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_5_15_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_5_15_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_5_15_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_5_15_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_4_15_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( dummy_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_5_14_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_6_15_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_4_15_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( dummy_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_5_14_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_6_15_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_4_15_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( dummy_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_5_14_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_6_15_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_5_15_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_5_15_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_5_15_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_5_15_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_5_15_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_5_15_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_5_15_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_5_15_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_5_15_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_5_15_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_5_15_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_5_15_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_4_15_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( dummy_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_5_14_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_6_15_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_4_15_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( dummy_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_5_14_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_6_15_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_4_15_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( dummy_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_5_14_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_6_15_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_5_15_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_5_15_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_5_15_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_5_15_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_5_15_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_5_15_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_5_15_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_5_15_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_5_15_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_5_15_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_5_15_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_5_15_out_S_noc3_yummy )
);


tile
tile111 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[111] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd15),
    .default_coreid_y           (8'd6),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd111)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[111]   )
    ,.unavailable_o       ( unavailable_o[111] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[111]   )
    ,.ipi_i               ( ipi_i[111]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[111*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile111_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile111_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_5_15_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( dummy_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_6_14_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_7_15_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_5_15_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( dummy_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_6_14_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_7_15_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_5_15_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( dummy_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_6_14_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_7_15_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_6_15_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_6_15_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_6_15_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_6_15_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_6_15_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_6_15_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_6_15_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_6_15_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_6_15_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_6_15_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_6_15_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_6_15_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_5_15_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( dummy_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_6_14_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_7_15_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_5_15_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( dummy_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_6_14_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_7_15_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_5_15_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( dummy_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_6_14_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_7_15_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_6_15_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_6_15_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_6_15_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_6_15_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_6_15_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_6_15_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_6_15_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_6_15_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_6_15_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_6_15_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_6_15_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_6_15_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_5_15_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( dummy_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_6_14_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_7_15_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_5_15_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( dummy_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_6_14_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_7_15_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_5_15_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( dummy_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_6_14_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_7_15_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_6_15_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_6_15_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_6_15_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_6_15_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_6_15_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_6_15_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_6_15_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_6_15_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_6_15_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_6_15_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_6_15_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_6_15_out_S_noc3_yummy )
);


tile
tile127 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[127] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd15),
    .default_coreid_y           (8'd7),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd127)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[127]   )
    ,.unavailable_o       ( unavailable_o[127] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[127]   )
    ,.ipi_i               ( ipi_i[127]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[127*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile127_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile127_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_6_15_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( dummy_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_7_14_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_8_15_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_6_15_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( dummy_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_7_14_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_8_15_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_6_15_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( dummy_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_7_14_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_8_15_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_7_15_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_7_15_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_7_15_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_7_15_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_7_15_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_7_15_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_7_15_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_7_15_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_7_15_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_7_15_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_7_15_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_7_15_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_6_15_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( dummy_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_7_14_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_8_15_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_6_15_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( dummy_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_7_14_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_8_15_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_6_15_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( dummy_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_7_14_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_8_15_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_7_15_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_7_15_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_7_15_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_7_15_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_7_15_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_7_15_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_7_15_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_7_15_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_7_15_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_7_15_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_7_15_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_7_15_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_6_15_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( dummy_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_7_14_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_8_15_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_6_15_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( dummy_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_7_14_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_8_15_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_6_15_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( dummy_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_7_14_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_8_15_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_7_15_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_7_15_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_7_15_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_7_15_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_7_15_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_7_15_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_7_15_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_7_15_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_7_15_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_7_15_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_7_15_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_7_15_out_S_noc3_yummy )
);


tile
tile143 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[143] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd15),
    .default_coreid_y           (8'd8),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd143)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[143]   )
    ,.unavailable_o       ( unavailable_o[143] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[143]   )
    ,.ipi_i               ( ipi_i[143]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[143*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile143_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile143_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_7_15_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( dummy_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_8_14_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_9_15_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_7_15_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( dummy_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_8_14_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_9_15_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_7_15_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( dummy_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_8_14_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_9_15_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_8_15_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_8_15_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_8_15_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_8_15_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_8_15_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_8_15_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_8_15_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_8_15_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_8_15_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_8_15_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_8_15_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_8_15_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_7_15_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( dummy_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_8_14_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_9_15_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_7_15_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( dummy_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_8_14_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_9_15_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_7_15_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( dummy_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_8_14_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_9_15_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_8_15_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_8_15_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_8_15_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_8_15_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_8_15_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_8_15_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_8_15_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_8_15_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_8_15_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_8_15_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_8_15_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_8_15_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_7_15_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( dummy_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_8_14_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_9_15_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_7_15_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( dummy_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_8_14_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_9_15_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_7_15_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( dummy_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_8_14_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_9_15_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_8_15_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_8_15_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_8_15_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_8_15_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_8_15_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_8_15_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_8_15_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_8_15_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_8_15_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_8_15_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_8_15_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_8_15_out_S_noc3_yummy )
);


tile
tile159 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[159] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd15),
    .default_coreid_y           (8'd9),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd159)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[159]   )
    ,.unavailable_o       ( unavailable_o[159] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[159]   )
    ,.ipi_i               ( ipi_i[159]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[159*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile159_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile159_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_8_15_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( dummy_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_9_14_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_10_15_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_8_15_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( dummy_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_9_14_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_10_15_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_8_15_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( dummy_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_9_14_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_10_15_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_9_15_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_9_15_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_9_15_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_9_15_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_9_15_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_9_15_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_9_15_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_9_15_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_9_15_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_9_15_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_9_15_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_9_15_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_8_15_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( dummy_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_9_14_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_10_15_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_8_15_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( dummy_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_9_14_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_10_15_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_8_15_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( dummy_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_9_14_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_10_15_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_9_15_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_9_15_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_9_15_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_9_15_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_9_15_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_9_15_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_9_15_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_9_15_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_9_15_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_9_15_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_9_15_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_9_15_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_8_15_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( dummy_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_9_14_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_10_15_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_8_15_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( dummy_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_9_14_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_10_15_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_8_15_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( dummy_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_9_14_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_10_15_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_9_15_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_9_15_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_9_15_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_9_15_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_9_15_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_9_15_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_9_15_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_9_15_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_9_15_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_9_15_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_9_15_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_9_15_out_S_noc3_yummy )
);


tile
tile175 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[175] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd15),
    .default_coreid_y           (8'd10),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd175)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[175]   )
    ,.unavailable_o       ( unavailable_o[175] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[175]   )
    ,.ipi_i               ( ipi_i[175]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[175*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile175_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile175_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_9_15_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( dummy_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_10_14_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_11_15_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_9_15_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( dummy_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_10_14_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_11_15_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_9_15_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( dummy_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_10_14_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_11_15_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_10_15_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_10_15_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_10_15_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_10_15_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_10_15_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_10_15_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_10_15_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_10_15_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_10_15_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_10_15_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_10_15_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_10_15_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_9_15_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( dummy_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_10_14_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_11_15_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_9_15_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( dummy_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_10_14_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_11_15_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_9_15_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( dummy_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_10_14_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_11_15_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_10_15_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_10_15_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_10_15_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_10_15_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_10_15_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_10_15_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_10_15_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_10_15_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_10_15_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_10_15_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_10_15_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_10_15_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_9_15_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( dummy_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_10_14_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_11_15_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_9_15_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( dummy_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_10_14_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_11_15_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_9_15_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( dummy_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_10_14_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_11_15_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_10_15_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_10_15_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_10_15_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_10_15_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_10_15_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_10_15_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_10_15_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_10_15_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_10_15_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_10_15_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_10_15_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_10_15_out_S_noc3_yummy )
);


tile
tile191 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[191] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd15),
    .default_coreid_y           (8'd11),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd191)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[191]   )
    ,.unavailable_o       ( unavailable_o[191] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[191]   )
    ,.ipi_i               ( ipi_i[191]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[191*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile191_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile191_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_10_15_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( dummy_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_11_14_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_12_15_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_10_15_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( dummy_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_11_14_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_12_15_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_10_15_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( dummy_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_11_14_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_12_15_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_11_15_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_11_15_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_11_15_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_11_15_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_11_15_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_11_15_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_11_15_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_11_15_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_11_15_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_11_15_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_11_15_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_11_15_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_10_15_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( dummy_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_11_14_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_12_15_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_10_15_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( dummy_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_11_14_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_12_15_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_10_15_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( dummy_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_11_14_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_12_15_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_11_15_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_11_15_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_11_15_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_11_15_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_11_15_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_11_15_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_11_15_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_11_15_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_11_15_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_11_15_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_11_15_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_11_15_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_10_15_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( dummy_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_11_14_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_12_15_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_10_15_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( dummy_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_11_14_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_12_15_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_10_15_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( dummy_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_11_14_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_12_15_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_11_15_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_11_15_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_11_15_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_11_15_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_11_15_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_11_15_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_11_15_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_11_15_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_11_15_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_11_15_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_11_15_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_11_15_out_S_noc3_yummy )
);


tile
tile207 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[207] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd15),
    .default_coreid_y           (8'd12),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd207)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[207]   )
    ,.unavailable_o       ( unavailable_o[207] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[207]   )
    ,.ipi_i               ( ipi_i[207]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[207*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile207_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile207_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_11_15_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( dummy_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_12_14_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_13_15_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_11_15_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( dummy_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_12_14_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_13_15_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_11_15_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( dummy_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_12_14_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_13_15_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_12_15_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_12_15_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_12_15_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_12_15_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_12_15_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_12_15_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_12_15_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_12_15_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_12_15_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_12_15_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_12_15_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_12_15_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_11_15_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( dummy_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_12_14_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_13_15_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_11_15_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( dummy_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_12_14_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_13_15_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_11_15_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( dummy_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_12_14_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_13_15_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_12_15_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_12_15_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_12_15_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_12_15_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_12_15_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_12_15_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_12_15_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_12_15_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_12_15_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_12_15_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_12_15_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_12_15_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_11_15_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( dummy_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_12_14_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_13_15_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_11_15_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( dummy_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_12_14_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_13_15_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_11_15_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( dummy_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_12_14_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_13_15_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_12_15_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_12_15_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_12_15_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_12_15_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_12_15_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_12_15_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_12_15_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_12_15_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_12_15_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_12_15_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_12_15_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_12_15_out_S_noc3_yummy )
);


tile
tile223 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[223] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd15),
    .default_coreid_y           (8'd13),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd223)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[223]   )
    ,.unavailable_o       ( unavailable_o[223] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[223]   )
    ,.ipi_i               ( ipi_i[223]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[223*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile223_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile223_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_12_15_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( dummy_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_13_14_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_14_15_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_12_15_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( dummy_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_13_14_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_14_15_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_12_15_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( dummy_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_13_14_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_14_15_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_13_15_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_13_15_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_13_15_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_13_15_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_13_15_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_13_15_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_13_15_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_13_15_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_13_15_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_13_15_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_13_15_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_13_15_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_12_15_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( dummy_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_13_14_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_14_15_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_12_15_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( dummy_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_13_14_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_14_15_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_12_15_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( dummy_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_13_14_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_14_15_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_13_15_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_13_15_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_13_15_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_13_15_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_13_15_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_13_15_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_13_15_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_13_15_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_13_15_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_13_15_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_13_15_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_13_15_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_12_15_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( dummy_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_13_14_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_14_15_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_12_15_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( dummy_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_13_14_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_14_15_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_12_15_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( dummy_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_13_14_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_14_15_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_13_15_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_13_15_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_13_15_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_13_15_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_13_15_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_13_15_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_13_15_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_13_15_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_13_15_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_13_15_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_13_15_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_13_15_out_S_noc3_yummy )
);


tile
tile239 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[239] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd15),
    .default_coreid_y           (8'd14),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd239)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[239]   )
    ,.unavailable_o       ( unavailable_o[239] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[239]   )
    ,.ipi_i               ( ipi_i[239]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[239*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile239_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile239_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_13_15_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( dummy_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_14_14_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( tile_15_15_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_13_15_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( dummy_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_14_14_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( tile_15_15_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_13_15_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( dummy_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_14_14_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( tile_15_15_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_14_15_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_14_15_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_14_15_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_14_15_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_14_15_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_14_15_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_14_15_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_14_15_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_14_15_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_14_15_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_14_15_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_14_15_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_13_15_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( dummy_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_14_14_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( tile_15_15_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_13_15_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( dummy_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_14_14_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( tile_15_15_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_13_15_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( dummy_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_14_14_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( tile_15_15_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_14_15_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_14_15_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_14_15_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_14_15_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_14_15_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_14_15_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_14_15_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_14_15_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_14_15_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_14_15_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_14_15_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_14_15_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_13_15_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( dummy_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_14_14_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( tile_15_15_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_13_15_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( dummy_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_14_14_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( tile_15_15_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_13_15_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( dummy_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_14_14_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( tile_15_15_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_14_15_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_14_15_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_14_15_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_14_15_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_14_15_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_14_15_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_14_15_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_14_15_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_14_15_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_14_15_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_14_15_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_14_15_out_S_noc3_yummy )
);


tile
tile255 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (/* ctap_clk_en_inter[255] always one */ 1'b1 && clk_en_inter),
    .default_chipid             (14'b0),    // the first chip
    .default_coreid_x           (8'd15),
    .default_coreid_y           (8'd15),
    .default_total_num_tiles    (default_total_num_tiles      ),
    .flat_tileid                (`JTAG_FLATID_WIDTH'd255)
`ifdef PITON_RV64_PLATFORM
`ifdef PITON_RV64_DEBUGUNIT
    ,.debug_req_i         ( debug_req_i[255]   )
    ,.unavailable_o       ( unavailable_o[255] )
`endif // ifdef PITON_RV64_DEBUGUNIT
`ifdef PITON_RV64_CLINT
    ,.timer_irq_i         ( timer_irq_i[255]   )
    ,.ipi_i               ( ipi_i[255]         )
`endif // ifdef PITON_RV64_CLINT
`ifdef PITON_RV64_PLIC
    ,.irq_i               ( irq_i[255*2 +: 2]  )
`endif // ifdef PITON_RV64_PLIC
`endif // ifdef PITON_RV64_PLATFORM
    ,
    // ucb from tiles to jtag
    .tile_jtag_ucb_val   ( tile255_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile255_jtag_ucb_data     ),
    // ucb from jtag to tiles
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),

    .dyn0_dataIn_N       ( tile_14_15_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( dummy_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( tile_15_14_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( dummy_out_N_noc1_data   ),
    .dyn0_validIn_N      ( tile_14_15_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( dummy_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( tile_15_14_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( dummy_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( tile_14_15_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( dummy_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( tile_15_14_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( dummy_out_N_noc1_yummy  ),

    .dyn0_dNo            ( tile_15_15_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_15_15_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_15_15_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_15_15_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_15_15_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_15_15_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_15_15_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_15_15_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_15_15_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_15_15_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_15_15_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_15_15_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( tile_14_15_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( dummy_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( tile_15_14_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( dummy_out_N_noc2_data   ),
    .dyn1_validIn_N      ( tile_14_15_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( dummy_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( tile_15_14_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( dummy_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( tile_14_15_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( dummy_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( tile_15_14_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( dummy_out_N_noc2_yummy  ),

    .dyn1_dNo            ( tile_15_15_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_15_15_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_15_15_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_15_15_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_15_15_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_15_15_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_15_15_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_15_15_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_15_15_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_15_15_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_15_15_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_15_15_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( tile_14_15_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( dummy_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( tile_15_14_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( dummy_out_N_noc3_data   ),
    .dyn2_validIn_N      ( tile_14_15_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( dummy_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( tile_15_14_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( dummy_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( tile_14_15_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( dummy_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( tile_15_14_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( dummy_out_N_noc3_yummy  ),

    .dyn2_dNo            ( tile_15_15_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_15_15_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_15_15_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_15_15_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_15_15_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_15_15_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_15_15_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_15_15_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_15_15_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_15_15_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_15_15_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_15_15_out_S_noc3_yummy )
);


endmodule

`endif
